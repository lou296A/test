

    module v_ROM1_462(q, a, clk);
    output reg [0:0] q;
    input [11:0] a;
    reg [0:0] rom [4095:0];
    always @(posedge clk) q <= rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end
    begin
        rom[0] = 0;
rom[1] = 1;
rom[2] = 0;
rom[3] = 0;
rom[4] = 0;
rom[5] = 1;
rom[6] = 0;
rom[7] = 0;
rom[8] = 0;
rom[9] = 1;
rom[10] = 1;
rom[11] = 1;
rom[12] = 0;
rom[13] = 0;
rom[14] = 1;
rom[15] = 0;
rom[16] = 0;
rom[17] = 0;
rom[18] = 0;
rom[19] = 0;
rom[20] = 0;
rom[21] = 1;
rom[22] = 1;
rom[23] = 1;
rom[24] = 1;
rom[25] = 0;
rom[26] = 0;
rom[27] = 0;
rom[28] = 0;
rom[29] = 0;
rom[30] = 0;
rom[31] = 1;
rom[32] = 1;
rom[33] = 1;
rom[34] = 1;
rom[35] = 1;
rom[36] = 1;
rom[37] = 1;
rom[38] = 1;
rom[39] = 1;
rom[40] = 1;
rom[41] = 1;
rom[42] = 1;
rom[43] = 1;
rom[44] = 1;
rom[45] = 1;
rom[46] = 1;
rom[47] = 1;
rom[48] = 1;
rom[49] = 1;
rom[50] = 1;
rom[51] = 1;
rom[52] = 1;
rom[53] = 1;
rom[54] = 1;
rom[55] = 1;
rom[56] = 1;
rom[57] = 1;
rom[58] = 1;
rom[59] = 1;
rom[60] = 1;
rom[61] = 1;
rom[62] = 1;
rom[63] = 1;
rom[64] = 1;
rom[65] = 1;
rom[66] = 1;
rom[67] = 1;
rom[68] = 1;
rom[69] = 1;
rom[70] = 1;
rom[71] = 1;
rom[72] = 1;
rom[73] = 1;
rom[74] = 1;
rom[75] = 1;
rom[76] = 1;
rom[77] = 1;
rom[78] = 1;
rom[79] = 1;
rom[80] = 1;
rom[81] = 1;
rom[82] = 1;
rom[83] = 1;
rom[84] = 1;
rom[85] = 1;
rom[86] = 1;
rom[87] = 1;
rom[88] = 1;
rom[89] = 1;
rom[90] = 1;
rom[91] = 1;
rom[92] = 1;
rom[93] = 1;
rom[94] = 1;
rom[95] = 1;
    end
     

    module v_RAM0_1680(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        ram[0] = 8192;
ram[1] = 838;
ram[2] = 1862;
ram[3] = 32769;
ram[4] = 1862;
ram[5] = 32769;
ram[6] = 322;
ram[7] = 28672;
ram[2036] = 50786;
ram[2037] = 205;
ram[2038] = 3281;
ram[2039] = 12997;
ram[2040] = 3797;
ram[2041] = 35840;
ram[2042] = 15561;
ram[2043] = 3285;
ram[2044] = 717;
ram[2045] = 3793;
ram[2046] = 50688;
    end
    endmodule

    

    module v_data_ram_1818(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        ram[0] = 15360;
ram[1] = 14336;
ram[2] = 12629;
ram[3] = 65535;
ram[4] = 8260;
ram[5] = 13312;
ram[6] = 85;
ram[7] = 0;
    end
    endmodule

    

    module v_RAM1_13398(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        ram[0] = 8192;
ram[1] = 722;
ram[2] = 3798;
ram[3] = 0;
ram[4] = 0;
ram[5] = 0;
ram[6] = 0;
ram[7] = 1742;
ram[8] = 32769;
ram[9] = 4099;
ram[10] = 28672;
ram[2036] = 50786;
ram[2037] = 205;
ram[2038] = 3281;
ram[2039] = 12997;
ram[2040] = 3797;
ram[2041] = 35840;
ram[2042] = 15561;
ram[2043] = 3285;
ram[2044] = 717;
ram[2045] = 3793;
ram[2046] = 50688;
    end
    endmodule

    
module main (
	clk,
	v_DIV_INST0_6905_out0,
	v_DIV_INST1_7011_out0,
	v_IR1_6873_out0,
	v_BYTE_RECEIVED_11192_out0,
	v_IR0_13305_out0,
	v_R13_375_out0,
	v_R11_398_out0,
	v_R00_3807_out0,
	v_R02_6966_out0,
	v_R12_10714_out0,
	v_R10_11216_out0,
	v_R03_13304_out0,
	v_R01_13752_out0,
	v_REGISTER_INUP16_384_out0,
	v_REGISTER_INUP0_12240_out0,
	v_REGISTER14_3201_out0,
	v_REGISTER15_8833_out0);
input clk;
input v_DIV_INST0_6905_out0;
input v_DIV_INST1_7011_out0;
output  [11:0] v_REGISTER14_3201_out0;
output  [11:0] v_REGISTER15_8833_out0;
output  [15:0] v_IR0_13305_out0;
output  [15:0] v_IR1_6873_out0;
output  [15:0] v_R00_3807_out0;
output  [15:0] v_R01_13752_out0;
output  [15:0] v_R02_6966_out0;
output  [15:0] v_R03_13304_out0;
output  [15:0] v_R10_11216_out0;
output  [15:0] v_R11_398_out0;
output  [15:0] v_R12_10714_out0;
output  [15:0] v_R13_375_out0;
output  [15:0] v_REGISTER_INUP0_12240_out0;
output  [15:0] v_REGISTER_INUP16_384_out0;
output  [7:0] v_BYTE_RECEIVED_11192_out0;
reg  [11:0] v_REG1_432_out0 = 12'h0;
reg  [11:0] v_REG1_433_out0 = 12'h0;
reg  [11:0] v_REG1_7134_out0 = 12'h0;
reg  [15:0] v_IHOLD_REGISTER_2013_out0 = 16'h0;
reg  [15:0] v_IHOLD_REGISTER_2014_out0 = 16'h0;
reg  [15:0] v_REG0_10912_out0 = 16'h0;
reg  [15:0] v_REG0_10913_out0 = 16'h0;
reg  [15:0] v_REG1_13338_out0 = 16'h0;
reg  [15:0] v_REG1_13339_out0 = 16'h0;
reg  [15:0] v_REG1_2314_out0 = 16'h0;
reg  [15:0] v_REG1_2315_out0 = 16'h0;
reg  [15:0] v_REG2_12251_out0 = 16'h0;
reg  [15:0] v_REG2_12252_out0 = 16'h0;
reg  [15:0] v_REG3_4747_out0 = 16'h0;
reg  [15:0] v_REG3_4748_out0 = 16'h0;
reg  [1:0] v_REG1_10368_out0 = 2'h0;
reg  [1:0] v_REG1_7031_out0 = 2'h0;
reg  [7:0] v_REG1_10546_out0 = 8'h0;
reg  [7:0] v_REG1_2677_out0 = 8'h0;
reg v_FF1_10325_out0 = 1'b0;
reg v_FF1_10326_out0 = 1'b0;
reg v_FF1_13511_out0 = 1'b0;
reg v_FF1_1955_out0 = 1'b0;
reg v_FF1_4717_out0 = 1'b0;
reg v_FF1_4718_out0 = 1'b0;
reg v_FF1_4719_out0 = 1'b0;
reg v_FF1_4720_out0 = 1'b0;
reg v_FF1_4721_out0 = 1'b0;
reg v_FF1_4722_out0 = 1'b0;
reg v_FF1_4723_out0 = 1'b0;
reg v_FF1_4724_out0 = 1'b0;
reg v_FF1_4725_out0 = 1'b0;
reg v_FF1_4726_out0 = 1'b0;
reg v_FF1_4727_out0 = 1'b0;
reg v_FF1_4728_out0 = 1'b0;
reg v_FF1_4729_out0 = 1'b0;
reg v_FF1_4730_out0 = 1'b0;
reg v_FF1_4731_out0 = 1'b0;
reg v_FF1_4732_out0 = 1'b0;
reg v_FF1_4841_out0 = 1'b0;
reg v_FF1_48_out0 = 1'b0;
reg v_FF1_49_out0 = 1'b0;
reg v_FF2_11062_out0 = 1'b0;
reg v_FF2_2833_out0 = 1'b0;
reg v_FF3_11046_out0 = 1'b0;
reg v_FF3_2016_out0 = 1'b0;
reg v_FF3_2017_out0 = 1'b0;
reg v_FF4_2106_out0 = 1'b0;
reg v_FF4_2107_out0 = 1'b0;
reg v_FF4_463_out0 = 1'b0;
reg v_FF5_7100_out0 = 1'b0;
reg v_FF6_112_out0 = 1'b0;
reg v_FF7_2670_out0 = 1'b0;
reg v_FF7_2671_out0 = 1'b0;
reg v_FF7_2672_out0 = 1'b0;
reg v_FF7_2673_out0 = 1'b0;
reg v_FF7_4781_out0 = 1'b0;
reg v_FF8_10849_out0 = 1'b0;
reg v_FF8_10850_out0 = 1'b0;
reg v_FF8_10851_out0 = 1'b0;
reg v_FF8_10852_out0 = 1'b0;
reg v_FF8_11222_out0 = 1'b0;
reg v_FF9_8805_out0 = 1'b0;
reg v_REG1_11130_out0 = 1'b0;
reg v_REG1_11131_out0 = 1'b0;
wire  [10:0] v_C1_606_out0;
wire  [10:0] v_C1_607_out0;
wire  [10:0] v_C_1807_out0;
wire  [10:0] v_C_1808_out0;
wire  [10:0] v_IN1_10992_out0;
wire  [10:0] v_IN1_10993_out0;
wire  [10:0] v_IN1_13711_out0;
wire  [10:0] v_IN1_13712_out0;
wire  [10:0] v_IN1_2189_out0;
wire  [10:0] v_IN1_2190_out0;
wire  [10:0] v_IN1_2848_out0;
wire  [10:0] v_IN1_2849_out0;
wire  [10:0] v_IN_13668_out0;
wire  [10:0] v_IN_13669_out0;
wire  [10:0] v_MUX1_2401_out0;
wire  [10:0] v_MUX1_2402_out0;
wire  [10:0] v_MUX1_7143_out0;
wire  [10:0] v_MUX1_7144_out0;
wire  [10:0] v_MUX1_7702_out0;
wire  [10:0] v_MUX1_7703_out0;
wire  [10:0] v_MUX2_188_out0;
wire  [10:0] v_MUX2_189_out0;
wire  [10:0] v_MUX3_13312_out0;
wire  [10:0] v_MUX3_13313_out0;
wire  [10:0] v_MUX4_552_out0;
wire  [10:0] v_MUX4_553_out0;
wire  [10:0] v_MUX5_13670_out0;
wire  [10:0] v_MUX5_13671_out0;
wire  [10:0] v_OP2_SIG11_14_out0;
wire  [10:0] v_OP2_SIG11_15_out0;
wire  [10:0] v_OP2_SIG11_4827_out0;
wire  [10:0] v_OP2_SIG11_4828_out0;
wire  [10:0] v_OP2_SIG_13314_out0;
wire  [10:0] v_OP2_SIG_13315_out0;
wire  [10:0] v_OP2_SIG_NEW_11190_out0;
wire  [10:0] v_OP2_SIG_NEW_11191_out0;
wire  [10:0] v_OP2_SIG_NEW_11218_out0;
wire  [10:0] v_OP2_SIG_NEW_11219_out0;
wire  [10:0] v_OUT1_1873_out0;
wire  [10:0] v_OUT1_1874_out0;
wire  [10:0] v_OUT1_1972_out0;
wire  [10:0] v_OUT1_1973_out0;
wire  [10:0] v_OUT1_3294_out0;
wire  [10:0] v_OUT1_3295_out0;
wire  [10:0] v_OUT1_3853_out0;
wire  [10:0] v_OUT1_3854_out0;
wire  [10:0] v_Q_10339_out0;
wire  [10:0] v_Q_10340_out0;
wire  [10:0] v_Q_10341_out0;
wire  [10:0] v_Q_10342_out0;
wire  [10:0] v_RD_SIG11_7132_out0;
wire  [10:0] v_RD_SIG11_7133_out0;
wire  [10:0] v_RD_SIG11_8854_out0;
wire  [10:0] v_RD_SIG11_8855_out0;
wire  [10:0] v_RD_SIG_109_out0;
wire  [10:0] v_RD_SIG_110_out0;
wire  [10:0] v_RD_SIG_NEW_10872_out0;
wire  [10:0] v_RD_SIG_NEW_10873_out0;
wire  [10:0] v_RD_SIG_NEW_8759_out0;
wire  [10:0] v_RD_SIG_NEW_8760_out0;
wire  [10:0] v_SEL2_13496_out0;
wire  [10:0] v_SEL2_13497_out0;
wire  [10:0] v_SHIFTED_SIG_10802_out0;
wire  [10:0] v_SHIFTED_SIG_10803_out0;
wire  [10:0] v_SHIFTED_SIG_13632_out0;
wire  [10:0] v_SHIFTED_SIG_13633_out0;
wire  [10:0] v_SIG_RD_11bit_3301_out0;
wire  [10:0] v_SIG_RD_11bit_3302_out0;
wire  [10:0] v_SIG_RM_11bit_6892_out0;
wire  [10:0] v_SIG_RM_11bit_6893_out0;
wire  [10:0] v_SIG_TO_SHIFT_10712_out0;
wire  [10:0] v_SIG_TO_SHIFT_10713_out0;
wire  [10:0] v_SIG_TO_SHIFT_5836_out0;
wire  [10:0] v_SIG_TO_SHIFT_5837_out0;
wire  [10:0] v__13310_out0;
wire  [10:0] v__13311_out0;
wire  [10:0] v__13484_out0;
wire  [10:0] v__13485_out0;
wire  [10:0] v__13761_out0;
wire  [10:0] v__13762_out0;
wire  [10:0] v__2026_out0;
wire  [10:0] v__2027_out0;
wire  [10:0] v__2028_out0;
wire  [10:0] v__2029_out0;
wire  [10:0] v__2030_out0;
wire  [10:0] v__2031_out0;
wire  [10:0] v__2032_out0;
wire  [10:0] v__2033_out0;
wire  [10:0] v__2034_out0;
wire  [10:0] v__2035_out0;
wire  [10:0] v__2036_out0;
wire  [10:0] v__2037_out0;
wire  [10:0] v__2038_out0;
wire  [10:0] v__2039_out0;
wire  [10:0] v__2040_out0;
wire  [10:0] v__2041_out0;
wire  [10:0] v__2042_out0;
wire  [10:0] v__2043_out0;
wire  [10:0] v__2044_out0;
wire  [10:0] v__2045_out0;
wire  [10:0] v__2046_out0;
wire  [10:0] v__2047_out0;
wire  [10:0] v__2048_out0;
wire  [10:0] v__2049_out0;
wire  [10:0] v__2050_out0;
wire  [10:0] v__2051_out0;
wire  [10:0] v__2052_out0;
wire  [10:0] v__2053_out0;
wire  [10:0] v__2054_out0;
wire  [10:0] v__2055_out0;
wire  [10:0] v__2191_out0;
wire  [10:0] v__2192_out0;
wire  [10:0] v__2771_out0;
wire  [10:0] v__2772_out0;
wire  [10:0] v__2834_out0;
wire  [10:0] v__2835_out0;
wire  [10:0] v__2836_out0;
wire  [10:0] v__2837_out0;
wire  [10:0] v__2971_out0;
wire  [10:0] v__2972_out0;
wire  [10:0] v__4591_out0;
wire  [10:0] v__4592_out0;
wire  [10:0] v__4733_out0;
wire  [10:0] v__4734_out0;
wire  [10:0] v__7714_out0;
wire  [10:0] v__7715_out0;
wire  [10:0] v_shifted1_2666_out0;
wire  [10:0] v_shifted1_2667_out0;
wire  [11:0] v_A1_11043_out0;
wire  [11:0] v_A1_7019_out0;
wire  [11:0] v_A1_7020_out0;
wire  [11:0] v_ADDER_IN_10995_out0;
wire  [11:0] v_ADDER_IN_10996_out0;
wire  [11:0] v_ADDRESS0_10982_out0;
wire  [11:0] v_ADDRESS1_2854_out0;
wire  [11:0] v_ADDRESS_4662_out0;
wire  [11:0] v_ADRESS0_11217_out0;
wire  [11:0] v_ADRESS1_1906_out0;
wire  [11:0] v_ADRESS_2339_out0;
wire  [11:0] v_ADRESS_2340_out0;
wire  [11:0] v_ADRESS_2542_out0;
wire  [11:0] v_ADRESS_2543_out0;
wire  [11:0] v_ADRESS_8683_out0;
wire  [11:0] v_ADRESS_ins0_11169_out0;
wire  [11:0] v_ADRESS_ins1_10617_out0;
wire  [11:0] v_A_10821_out0;
wire  [11:0] v_A_10822_out0;
wire  [11:0] v_C1_2426_out0;
wire  [11:0] v_C1_2427_out0;
wire  [11:0] v_C1_3210_out0;
wire  [11:0] v_C1_3211_out0;
wire  [11:0] v_C2_10761_out0;
wire  [11:0] v_C2_10762_out0;
wire  [11:0] v_C2_2413_out0;
wire  [11:0] v_EA_13516_out0;
wire  [11:0] v_EA_13517_out0;
wire  [11:0] v_JUMPADRESS_4745_out0;
wire  [11:0] v_JUMPADRESS_4746_out0;
wire  [11:0] v_JUMPADRESS_6964_out0;
wire  [11:0] v_JUMPADRESS_6965_out0;
wire  [11:0] v_MULTI_PRODUCT_7104_out0;
wire  [11:0] v_MULTI_PRODUCT_7105_out0;
wire  [11:0] v_MUX1_10773_out0;
wire  [11:0] v_MUX1_10774_out0;
wire  [11:0] v_MUX1_7097_out0;
wire  [11:0] v_MUX2_13656_out0;
wire  [11:0] v_MUX2_13657_out0;
wire  [11:0] v_MUX3_10330_out0;
wire  [11:0] v_MUX3_10331_out0;
wire  [11:0] v_MUX3_3225_out0;
wire  [11:0] v_MUX3_3226_out0;
wire  [11:0] v_MUX4_2658_out0;
wire  [11:0] v_MUX4_2659_out0;
wire  [11:0] v_MUX5_10845_out0;
wire  [11:0] v_MUX5_10846_out0;
wire  [11:0] v_MUX8_13785_out0;
wire  [11:0] v_MUX8_13786_out0;
wire  [11:0] v_NEXTADD_10526_out0;
wire  [11:0] v_NEXTADD_10527_out0;
wire  [11:0] v_NEXTADRESS_1803_out0;
wire  [11:0] v_NEXTADRESS_1804_out0;
wire  [11:0] v_NEXT_ADRESS_3243_out0;
wire  [11:0] v_NEXT_ADRESS_3244_out0;
wire  [11:0] v_NOUSED_13492_out0;
wire  [11:0] v_NOUSED_13493_out0;
wire  [11:0] v_PC_COUNTER_25_out0;
wire  [11:0] v_PC_COUNTER_26_out0;
wire  [11:0] v_PC_COUNTER_NEXT_7064_out0;
wire  [11:0] v_PC_COUNTER_NEXT_7065_out0;
wire  [11:0] v_RAMADDRMUX_10542_out0;
wire  [11:0] v_RAMADDRMUX_10543_out0;
wire  [11:0] v_RAMADDRMUX_2232_out0;
wire  [11:0] v_RAMADDRMUX_2233_out0;
wire  [11:0] v_RAMADDRMUX_7066_out0;
wire  [11:0] v_RAMADDRMUX_7067_out0;
wire  [11:0] v_RAMADDRMUX_92_out0;
wire  [11:0] v_RAMADDRMUX_93_out0;
wire  [11:0] v_RAM_ADDRESS_MUX_8803_out0;
wire  [11:0] v_RAM_ADDRESS_MUX_8804_out0;
wire  [11:0] v_RAM_ADDRES_MUX_13649_out0;
wire  [11:0] v_RAM_ADDRES_MUX_13650_out0;
wire  [11:0] v_REGISTER4_1705_out0;
wire  [11:0] v_REGISTER4_1706_out0;
wire  [11:0] v_REGISTER_13346_out0;
wire  [11:0] v_REGISTER_13347_out0;
wire  [11:0] v_REGISTER_216_out0;
wire  [11:0] v_REGISTER_217_out0;
wire  [11:0] v_SEL7_4850_out0;
wire  [11:0] v_SEL7_4851_out0;
wire  [11:0] v_SEL8_10686_out0;
wire  [11:0] v_SEL8_10687_out0;
wire  [11:0] v__10370_out0;
wire  [11:0] v__10371_out0;
wire  [11:0] v__10783_out0;
wire  [11:0] v__10784_out0;
wire  [11:0] v__107_out0;
wire  [11:0] v__108_out0;
wire  [11:0] v__11137_out0;
wire  [11:0] v__11138_out0;
wire  [11:0] v__11139_out0;
wire  [11:0] v__11140_out0;
wire  [11:0] v__13291_out1;
wire  [11:0] v__13292_out1;
wire  [11:0] v__224_out0;
wire  [11:0] v__225_out0;
wire  [11:0] v__2411_out0;
wire  [11:0] v__2412_out0;
wire  [11:0] v__2439_out0;
wire  [11:0] v__2440_out0;
wire  [11:0] v__2793_out0;
wire  [11:0] v__2794_out0;
wire  [11:0] v__2795_out0;
wire  [11:0] v__2796_out0;
wire  [11:0] v__2797_out0;
wire  [11:0] v__2798_out0;
wire  [11:0] v__2799_out0;
wire  [11:0] v__2800_out0;
wire  [11:0] v__2801_out0;
wire  [11:0] v__2802_out0;
wire  [11:0] v__2803_out0;
wire  [11:0] v__2804_out0;
wire  [11:0] v__2805_out0;
wire  [11:0] v__2806_out0;
wire  [11:0] v__2807_out0;
wire  [11:0] v__2808_out0;
wire  [11:0] v__2809_out0;
wire  [11:0] v__2810_out0;
wire  [11:0] v__2811_out0;
wire  [11:0] v__2812_out0;
wire  [11:0] v__2813_out0;
wire  [11:0] v__2814_out0;
wire  [11:0] v__2815_out0;
wire  [11:0] v__2816_out0;
wire  [11:0] v__2817_out0;
wire  [11:0] v__2818_out0;
wire  [11:0] v__2819_out0;
wire  [11:0] v__2820_out0;
wire  [11:0] v__2821_out0;
wire  [11:0] v__2822_out0;
wire  [11:0] v__3035_out0;
wire  [11:0] v__3036_out0;
wire  [11:0] v__4488_out1;
wire  [11:0] v__4489_out1;
wire  [11:0] v__4585_out1;
wire  [11:0] v__4586_out1;
wire  [11:0] v__5846_out0;
wire  [11:0] v__5847_out0;
wire  [11:0] v__7116_out0;
wire  [11:0] v__7117_out0;
wire  [12:0] v__164_out0;
wire  [12:0] v__165_out0;
wire  [12:0] v__1825_out0;
wire  [12:0] v__1826_out0;
wire  [12:0] v__1827_out0;
wire  [12:0] v__1828_out0;
wire  [12:0] v__1829_out0;
wire  [12:0] v__1830_out0;
wire  [12:0] v__1831_out0;
wire  [12:0] v__1832_out0;
wire  [12:0] v__1833_out0;
wire  [12:0] v__1834_out0;
wire  [12:0] v__1835_out0;
wire  [12:0] v__1836_out0;
wire  [12:0] v__1837_out0;
wire  [12:0] v__1838_out0;
wire  [12:0] v__1839_out0;
wire  [12:0] v__1840_out0;
wire  [12:0] v__1841_out0;
wire  [12:0] v__1842_out0;
wire  [12:0] v__1843_out0;
wire  [12:0] v__1844_out0;
wire  [12:0] v__1845_out0;
wire  [12:0] v__1846_out0;
wire  [12:0] v__1847_out0;
wire  [12:0] v__1848_out0;
wire  [12:0] v__1849_out0;
wire  [12:0] v__1850_out0;
wire  [12:0] v__1851_out0;
wire  [12:0] v__1852_out0;
wire  [12:0] v__1853_out0;
wire  [12:0] v__1854_out0;
wire  [12:0] v__3192_out0;
wire  [12:0] v__3193_out0;
wire  [12:0] v__3194_out0;
wire  [12:0] v__3195_out0;
wire  [12:0] v__5851_out0;
wire  [12:0] v__5852_out0;
wire  [12:0] v__9802_out0;
wire  [12:0] v__9803_out0;
wire  [13:0] v__10767_out0;
wire  [13:0] v__10768_out0;
wire  [13:0] v__11049_out0;
wire  [13:0] v__11050_out0;
wire  [13:0] v__11055_out0;
wire  [13:0] v__11056_out0;
wire  [13:0] v__173_out0;
wire  [13:0] v__174_out0;
wire  [13:0] v__175_out0;
wire  [13:0] v__176_out0;
wire  [13:0] v__4483_out1;
wire  [13:0] v__4484_out1;
wire  [13:0] v__4549_out0;
wire  [13:0] v__4550_out0;
wire  [13:0] v__4551_out0;
wire  [13:0] v__4552_out0;
wire  [13:0] v__4553_out0;
wire  [13:0] v__4554_out0;
wire  [13:0] v__4555_out0;
wire  [13:0] v__4556_out0;
wire  [13:0] v__4557_out0;
wire  [13:0] v__4558_out0;
wire  [13:0] v__4559_out0;
wire  [13:0] v__4560_out0;
wire  [13:0] v__4561_out0;
wire  [13:0] v__4562_out0;
wire  [13:0] v__4563_out0;
wire  [13:0] v__4564_out0;
wire  [13:0] v__4565_out0;
wire  [13:0] v__4566_out0;
wire  [13:0] v__4567_out0;
wire  [13:0] v__4568_out0;
wire  [13:0] v__4569_out0;
wire  [13:0] v__4570_out0;
wire  [13:0] v__4571_out0;
wire  [13:0] v__4572_out0;
wire  [13:0] v__4573_out0;
wire  [13:0] v__4574_out0;
wire  [13:0] v__4575_out0;
wire  [13:0] v__4576_out0;
wire  [13:0] v__4577_out0;
wire  [13:0] v__4578_out0;
wire  [13:0] v__4816_out1;
wire  [13:0] v__4817_out1;
wire  [13:0] v__538_out0;
wire  [13:0] v__539_out0;
wire  [13:0] v__627_out1;
wire  [13:0] v__628_out1;
wire  [14:0] v_CIN_2356_out0;
wire  [14:0] v_CIN_2371_out0;
wire  [14:0] v_REST_162_out0;
wire  [14:0] v_REST_163_out0;
wire  [14:0] v__10354_out0;
wire  [14:0] v__10355_out0;
wire  [14:0] v__10455_out0;
wire  [14:0] v__10456_out0;
wire  [14:0] v__10457_out0;
wire  [14:0] v__10458_out0;
wire  [14:0] v__10651_out0;
wire  [14:0] v__10652_out0;
wire  [14:0] v__10653_out0;
wire  [14:0] v__10654_out0;
wire  [14:0] v__10655_out0;
wire  [14:0] v__10656_out0;
wire  [14:0] v__10657_out0;
wire  [14:0] v__10658_out0;
wire  [14:0] v__10659_out0;
wire  [14:0] v__10660_out0;
wire  [14:0] v__10661_out0;
wire  [14:0] v__10662_out0;
wire  [14:0] v__10663_out0;
wire  [14:0] v__10664_out0;
wire  [14:0] v__10665_out0;
wire  [14:0] v__10666_out0;
wire  [14:0] v__10667_out0;
wire  [14:0] v__10668_out0;
wire  [14:0] v__10669_out0;
wire  [14:0] v__10670_out0;
wire  [14:0] v__10671_out0;
wire  [14:0] v__10672_out0;
wire  [14:0] v__10673_out0;
wire  [14:0] v__10674_out0;
wire  [14:0] v__10675_out0;
wire  [14:0] v__10676_out0;
wire  [14:0] v__10677_out0;
wire  [14:0] v__10678_out0;
wire  [14:0] v__10679_out0;
wire  [14:0] v__10680_out0;
wire  [14:0] v__10910_out1;
wire  [14:0] v__10911_out1;
wire  [14:0] v__11231_out0;
wire  [14:0] v__11232_out0;
wire  [14:0] v__11294_out0;
wire  [14:0] v__11295_out0;
wire  [14:0] v__13709_out0;
wire  [14:0] v__13710_out0;
wire  [14:0] v__2223_out0;
wire  [14:0] v__2224_out0;
wire  [14:0] v__2889_out1;
wire  [14:0] v__2890_out1;
wire  [14:0] v__2984_out1;
wire  [14:0] v__2985_out1;
wire  [14:0] v__4831_out0;
wire  [14:0] v__4832_out0;
wire  [14:0] v__4856_out1;
wire  [14:0] v__4857_out1;
wire  [15:0] v_16BIT_WORD_ANSWER_8821_out0;
wire  [15:0] v_16BIT_WORD_ANSWER_8822_out0;
wire  [15:0] v_A1_3174_out0;
wire  [15:0] v_A1_3175_out0;
wire  [15:0] v_A1_3855_out0;
wire  [15:0] v_A1_3856_out0;
wire  [15:0] v_A4_11227_out0;
wire  [15:0] v_A4_11228_out0;
wire  [15:0] v_A5_1901_out0;
wire  [15:0] v_A5_1902_out0;
wire  [15:0] v_A6_10463_out0;
wire  [15:0] v_A6_10464_out0;
wire  [15:0] v_A8_11155_out0;
wire  [15:0] v_A8_11156_out0;
wire  [15:0] v_ADDER_IN_8744_out0;
wire  [15:0] v_ADDER_IN_8745_out0;
wire  [15:0] v_ADDER_IN_8746_out0;
wire  [15:0] v_ADDER_IN_8747_out0;
wire  [15:0] v_ALUOUT_10528_out0;
wire  [15:0] v_ALUOUT_10529_out0;
wire  [15:0] v_ALUOUT_11053_out0;
wire  [15:0] v_ALUOUT_11054_out0;
wire  [15:0] v_ALUOUT_4494_out0;
wire  [15:0] v_ALUOUT_4495_out0;
wire  [15:0] v_ALUOUT_4607_out0;
wire  [15:0] v_ALUOUT_4608_out0;
wire  [15:0] v_ALUOUT_8856_out0;
wire  [15:0] v_ALUOUT_8857_out0;
wire  [15:0] v_ANDOUT_630_out0;
wire  [15:0] v_ANDOUT_631_out0;
wire  [15:0] v_ANDOUT_632_out0;
wire  [15:0] v_ANDOUT_633_out0;
wire  [15:0] v_A_10274_out0;
wire  [15:0] v_A_10275_out0;
wire  [15:0] v_A_10276_out0;
wire  [15:0] v_A_10277_out0;
wire  [15:0] v_A_11250_out0;
wire  [15:0] v_A_11251_out0;
wire  [15:0] v_A_11252_out0;
wire  [15:0] v_A_11253_out0;
wire  [15:0] v_B_3350_out0;
wire  [15:0] v_B_3352_out0;
wire  [15:0] v_C11_4539_out0;
wire  [15:0] v_C11_4540_out0;
wire  [15:0] v_C13_2185_out0;
wire  [15:0] v_C13_2186_out0;
wire  [15:0] v_C15_1730_out0;
wire  [15:0] v_C15_1731_out0;
wire  [15:0] v_C5_2688_out0;
wire  [15:0] v_C5_2689_out0;
wire  [15:0] v_C7_1865_out0;
wire  [15:0] v_C7_1866_out0;
wire  [15:0] v_CIN_2355_out0;
wire  [15:0] v_CIN_2357_out0;
wire  [15:0] v_CIN_2358_out0;
wire  [15:0] v_CIN_2359_out0;
wire  [15:0] v_CIN_2360_out0;
wire  [15:0] v_CIN_2361_out0;
wire  [15:0] v_CIN_2362_out0;
wire  [15:0] v_CIN_2363_out0;
wire  [15:0] v_CIN_2364_out0;
wire  [15:0] v_CIN_2365_out0;
wire  [15:0] v_CIN_2366_out0;
wire  [15:0] v_CIN_2367_out0;
wire  [15:0] v_CIN_2368_out0;
wire  [15:0] v_CIN_2369_out0;
wire  [15:0] v_CIN_2370_out0;
wire  [15:0] v_CIN_2372_out0;
wire  [15:0] v_CIN_2373_out0;
wire  [15:0] v_CIN_2374_out0;
wire  [15:0] v_CIN_2375_out0;
wire  [15:0] v_CIN_2376_out0;
wire  [15:0] v_CIN_2377_out0;
wire  [15:0] v_CIN_2378_out0;
wire  [15:0] v_CIN_2379_out0;
wire  [15:0] v_CIN_2380_out0;
wire  [15:0] v_CIN_2381_out0;
wire  [15:0] v_CIN_2382_out0;
wire  [15:0] v_CIN_2383_out0;
wire  [15:0] v_CIN_2384_out0;
wire  [15:0] v_COUT_10916_out0;
wire  [15:0] v_COUT_10917_out0;
wire  [15:0] v_COUT_10918_out0;
wire  [15:0] v_COUT_10919_out0;
wire  [15:0] v_COUT_10920_out0;
wire  [15:0] v_COUT_10921_out0;
wire  [15:0] v_COUT_10922_out0;
wire  [15:0] v_COUT_10923_out0;
wire  [15:0] v_COUT_10924_out0;
wire  [15:0] v_COUT_10925_out0;
wire  [15:0] v_COUT_10926_out0;
wire  [15:0] v_COUT_10927_out0;
wire  [15:0] v_COUT_10928_out0;
wire  [15:0] v_COUT_10929_out0;
wire  [15:0] v_COUT_10930_out0;
wire  [15:0] v_COUT_10931_out0;
wire  [15:0] v_COUT_10932_out0;
wire  [15:0] v_COUT_10933_out0;
wire  [15:0] v_COUT_10934_out0;
wire  [15:0] v_COUT_10935_out0;
wire  [15:0] v_COUT_10936_out0;
wire  [15:0] v_COUT_10937_out0;
wire  [15:0] v_COUT_10938_out0;
wire  [15:0] v_COUT_10939_out0;
wire  [15:0] v_COUT_10940_out0;
wire  [15:0] v_COUT_10941_out0;
wire  [15:0] v_COUT_10942_out0;
wire  [15:0] v_COUT_10943_out0;
wire  [15:0] v_COUT_10944_out0;
wire  [15:0] v_COUT_10945_out0;
wire  [15:0] v_DATA0_13293_out0;
wire  [15:0] v_DATA0_4737_out0;
wire  [15:0] v_DATA1_1974_out0;
wire  [15:0] v_DATA1_603_out0;
wire  [15:0] v_DATA_10445_out0;
wire  [15:0] v_DATA_2469_out0;
wire  [15:0] v_DATA_IN_10552_out0;
wire  [15:0] v_DATA_IN_10553_out0;
wire  [15:0] v_DATA_OUT_1135_out0;
wire  [15:0] v_DATA_RAM_IN0_284_out0;
wire  [15:0] v_DATA_RAM_IN1_4779_out0;
wire  [15:0] v_DATA_RAM_IN_558_out0;
wire  [15:0] v_DATA_RAM_IN_559_out0;
wire  [15:0] v_DATA_to_transmit_4546_out0;
wire  [15:0] v_DFQDF_3025_out0;
wire  [15:0] v_DFQDF_3026_out0;
wire  [15:0] v_DIN3_10310_out0;
wire  [15:0] v_DIN3_10311_out0;
wire  [15:0] v_DIN_2266_out0;
wire  [15:0] v_DIN_2267_out0;
wire  [15:0] v_DIN_9798_out0;
wire  [15:0] v_DIN_9799_out0;
wire  [15:0] v_DOUT1_1207_out0;
wire  [15:0] v_DOUT1_1208_out0;
wire  [15:0] v_DOUT2_1733_out0;
wire  [15:0] v_DOUT2_1734_out0;
wire  [15:0] v_FLOATING_REGISTER_IN_562_out0;
wire  [15:0] v_FLOATING_REGISTER_IN_563_out0;
wire  [15:0] v_IN_10403_out0;
wire  [15:0] v_IN_10404_out0;
wire  [15:0] v_IN_11258_out0;
wire  [15:0] v_IN_11259_out0;
wire  [15:0] v_IN_13306_out0;
wire  [15:0] v_IN_13307_out0;
wire  [15:0] v_IN_13548_out0;
wire  [15:0] v_IN_13549_out0;
wire  [15:0] v_IN_13788_out0;
wire  [15:0] v_IN_13789_out0;
wire  [15:0] v_IN_190_out0;
wire  [15:0] v_IN_191_out0;
wire  [15:0] v_IN_1964_out0;
wire  [15:0] v_IN_1965_out0;
wire  [15:0] v_IN_2350_out0;
wire  [15:0] v_IN_2351_out0;
wire  [15:0] v_IN_2664_out0;
wire  [15:0] v_IN_2665_out0;
wire  [15:0] v_IN_5796_out0;
wire  [15:0] v_IN_5797_out0;
wire  [15:0] v_IN_685_out0;
wire  [15:0] v_IN_686_out0;
wire  [15:0] v_IN_8838_out0;
wire  [15:0] v_IN_8839_out0;
wire  [15:0] v_IN_98_out0;
wire  [15:0] v_IN_99_out0;
wire  [15:0] v_IR_105_out0;
wire  [15:0] v_IR_106_out0;
wire  [15:0] v_IR_10816_out0;
wire  [15:0] v_IR_10817_out0;
wire  [15:0] v_IR_13480_out0;
wire  [15:0] v_IR_13481_out0;
wire  [15:0] v_IR_1871_out0;
wire  [15:0] v_IR_1872_out0;
wire  [15:0] v_IR_2826_out0;
wire  [15:0] v_IR_2827_out0;
wire  [15:0] v_IR_2901_out0;
wire  [15:0] v_IR_2902_out0;
wire  [15:0] v_IR_640_out0;
wire  [15:0] v_IR_641_out0;
wire  [15:0] v_IR_7112_out0;
wire  [15:0] v_IR_7113_out0;
wire  [15:0] v_IR_7706_out0;
wire  [15:0] v_IR_7707_out0;
wire  [15:0] v_KEXTEND_13329_out0;
wire  [15:0] v_KEXTEND_13330_out0;
wire  [15:0] v_LS_REGIN_3303_out0;
wire  [15:0] v_LS_REGIN_3304_out0;
wire  [15:0] v_MEM_RAM_434_out0;
wire  [15:0] v_MEM_RAM_435_out0;
wire  [15:0] v_MULTI_OUT_13607_out0;
wire  [15:0] v_MULTI_OUT_13608_out0;
wire  [15:0] v_MULTI_OUT_1669_out0;
wire  [15:0] v_MULTI_OUT_1670_out0;
wire  [15:0] v_MULTI_REGIN_2870_out0;
wire  [15:0] v_MULTI_REGIN_2871_out0;
wire  [15:0] v_MUX11_13745_out0;
wire  [15:0] v_MUX11_13746_out0;
wire  [15:0] v_MUX12_1714_out0;
wire  [15:0] v_MUX12_1715_out0;
wire  [15:0] v_MUX1_10443_out0;
wire  [15:0] v_MUX1_10444_out0;
wire  [15:0] v_MUX1_11141_out0;
wire  [15:0] v_MUX1_11142_out0;
wire  [15:0] v_MUX1_1735_out0;
wire  [15:0] v_MUX1_1736_out0;
wire  [15:0] v_MUX1_1883_out0;
wire  [15:0] v_MUX1_1884_out0;
wire  [15:0] v_MUX1_2532_out0;
wire  [15:0] v_MUX1_2533_out0;
wire  [15:0] v_MUX1_2717_out0;
wire  [15:0] v_MUX1_2718_out0;
wire  [15:0] v_MUX1_31_out0;
wire  [15:0] v_MUX1_32_out0;
wire  [15:0] v_MUX1_4844_out0;
wire  [15:0] v_MUX1_4845_out0;
wire  [15:0] v_MUX1_6_out0;
wire  [15:0] v_MUX1_7_out0;
wire  [15:0] v_MUX1_8813_out0;
wire  [15:0] v_MUX1_8814_out0;
wire  [15:0] v_MUX2_10841_out0;
wire  [15:0] v_MUX2_10842_out0;
wire  [15:0] v_MUX2_1181_out0;
wire  [15:0] v_MUX2_1182_out0;
wire  [15:0] v_MUX2_1199_out0;
wire  [15:0] v_MUX2_1200_out0;
wire  [15:0] v_MUX2_13319_out0;
wire  [15:0] v_MUX2_13320_out0;
wire  [15:0] v_MUX2_2337_out0;
wire  [15:0] v_MUX2_2338_out0;
wire  [15:0] v_MUX2_3202_out0;
wire  [15:0] v_MUX2_3203_out0;
wire  [15:0] v_MUX2_3255_out0;
wire  [15:0] v_MUX2_3256_out0;
wire  [15:0] v_MUX2_4612_out0;
wire  [15:0] v_MUX2_4613_out0;
wire  [15:0] v_MUX3_10787_out0;
wire  [15:0] v_MUX3_13335_out0;
wire  [15:0] v_MUX3_13336_out0;
wire  [15:0] v_MUX3_2058_out0;
wire  [15:0] v_MUX3_2059_out0;
wire  [15:0] v_MUX3_3041_out0;
wire  [15:0] v_MUX3_3042_out0;
wire  [15:0] v_MUX3_3133_out0;
wire  [15:0] v_MUX3_3134_out0;
wire  [15:0] v_MUX3_313_out0;
wire  [15:0] v_MUX3_314_out0;
wire  [15:0] v_MUX3_6864_out0;
wire  [15:0] v_MUX3_6865_out0;
wire  [15:0] v_MUX3_7075_out0;
wire  [15:0] v_MUX3_7076_out0;
wire  [15:0] v_MUX3_8669_out0;
wire  [15:0] v_MUX3_8670_out0;
wire  [15:0] v_MUX4_10524_out0;
wire  [15:0] v_MUX4_10525_out0;
wire  [15:0] v_MUX4_10_out0;
wire  [15:0] v_MUX4_11_out0;
wire  [15:0] v_MUX4_13498_out0;
wire  [15:0] v_MUX4_13499_out0;
wire  [15:0] v_MUX4_1698_out0;
wire  [15:0] v_MUX4_2229_out0;
wire  [15:0] v_MUX4_2230_out0;
wire  [15:0] v_MUX4_376_out0;
wire  [15:0] v_MUX4_377_out0;
wire  [15:0] v_MUX4_4579_out0;
wire  [15:0] v_MUX4_4580_out0;
wire  [15:0] v_MUX4_7023_out0;
wire  [15:0] v_MUX4_7024_out0;
wire  [15:0] v_MUX5_10605_out0;
wire  [15:0] v_MUX5_10606_out0;
wire  [15:0] v_MUX5_1185_out0;
wire  [15:0] v_MUX5_1186_out0;
wire  [15:0] v_MUX5_2595_out0;
wire  [15:0] v_MUX5_2596_out0;
wire  [15:0] v_MUX5_2606_out0;
wire  [15:0] v_MUX5_2607_out0;
wire  [15:0] v_MUX5_3305_out0;
wire  [15:0] v_MUX5_3306_out0;
wire  [15:0] v_MUX5_7017_out0;
wire  [15:0] v_MUX5_7018_out0;
wire  [15:0] v_MUX5_8840_out0;
wire  [15:0] v_MUX5_8841_out0;
wire  [15:0] v_MUX6_2341_out0;
wire  [15:0] v_MUX6_2342_out0;
wire  [15:0] v_MUX7_1165_out0;
wire  [15:0] v_MUX7_1166_out0;
wire  [15:0] v_MUX8_1907_out0;
wire  [15:0] v_MUX8_1908_out0;
wire  [15:0] v_M_REGIN_271_out0;
wire  [15:0] v_M_REGIN_272_out0;
wire  [15:0] v_OP1_2060_out0;
wire  [15:0] v_OP1_2061_out0;
wire  [15:0] v_OP1_2979_out0;
wire  [15:0] v_OP1_2980_out0;
wire  [15:0] v_OP1_3899_out0;
wire  [15:0] v_OP1_3900_out0;
wire  [15:0] v_OP2_10751_out0;
wire  [15:0] v_OP2_10752_out0;
wire  [15:0] v_OP2_11153_out0;
wire  [15:0] v_OP2_11154_out0;
wire  [15:0] v_OP2_2322_out0;
wire  [15:0] v_OP2_2323_out0;
wire  [15:0] v_OP2_2862_out0;
wire  [15:0] v_OP2_2863_out0;
wire  [15:0] v_OP2_3940_out0;
wire  [15:0] v_OP2_3941_out0;
wire  [15:0] v_OUT_10264_out0;
wire  [15:0] v_OUT_10265_out0;
wire  [15:0] v_OUT_11234_out0;
wire  [15:0] v_OUT_11235_out0;
wire  [15:0] v_OUT_1136_out0;
wire  [15:0] v_OUT_1137_out0;
wire  [15:0] v_OUT_12236_out0;
wire  [15:0] v_OUT_12237_out0;
wire  [15:0] v_OUT_2352_out0;
wire  [15:0] v_OUT_2353_out0;
wire  [15:0] v_OUT_2857_out0;
wire  [15:0] v_OUT_2858_out0;
wire  [15:0] v_OUT_460_out0;
wire  [15:0] v_OUT_461_out0;
wire  [15:0] v_OUT_7708_out0;
wire  [15:0] v_OUT_7709_out0;
wire  [15:0] v_OUT_7710_out0;
wire  [15:0] v_OUT_7711_out0;
wire  [15:0] v_OUT_8852_out0;
wire  [15:0] v_OUT_8853_out0;
wire  [15:0] v_R0TEST_3184_out0;
wire  [15:0] v_R0TEST_3185_out0;
wire  [15:0] v_R0TEST_7005_out0;
wire  [15:0] v_R0TEST_7006_out0;
wire  [15:0] v_R0_13295_out0;
wire  [15:0] v_R0_13296_out0;
wire  [15:0] v_R0_1688_out0;
wire  [15:0] v_R0_1689_out0;
wire  [15:0] v_R0_2537_out0;
wire  [15:0] v_R0_2538_out0;
wire  [15:0] v_R0_2850_out0;
wire  [15:0] v_R0_2851_out0;
wire  [15:0] v_R1TEST_10485_out0;
wire  [15:0] v_R1TEST_10486_out0;
wire  [15:0] v_R1TEST_10498_out0;
wire  [15:0] v_R1TEST_10499_out0;
wire  [15:0] v_R1_2056_out0;
wire  [15:0] v_R1_2057_out0;
wire  [15:0] v_R1_2630_out0;
wire  [15:0] v_R1_2631_out0;
wire  [15:0] v_R1_2723_out0;
wire  [15:0] v_R1_2724_out0;
wire  [15:0] v_R1_8761_out0;
wire  [15:0] v_R1_8762_out0;
wire  [15:0] v_R2TEST_10708_out0;
wire  [15:0] v_R2TEST_10709_out0;
wire  [15:0] v_R2TEST_10987_out0;
wire  [15:0] v_R2TEST_10988_out0;
wire  [15:0] v_R2_10556_out0;
wire  [15:0] v_R2_10557_out0;
wire  [15:0] v_R2_10904_out0;
wire  [15:0] v_R2_10905_out0;
wire  [15:0] v_R2_1726_out0;
wire  [15:0] v_R2_1727_out0;
wire  [15:0] v_R2_3043_out0;
wire  [15:0] v_R2_3044_out0;
wire  [15:0] v_R3TEST_117_out0;
wire  [15:0] v_R3TEST_118_out0;
wire  [15:0] v_R3TEST_2872_out0;
wire  [15:0] v_R3TEST_2873_out0;
wire  [15:0] v_R3_27_out0;
wire  [15:0] v_R3_28_out0;
wire  [15:0] v_R3_33_out0;
wire  [15:0] v_R3_34_out0;
wire  [15:0] v_R3_4652_out0;
wire  [15:0] v_R3_4653_out0;
wire  [15:0] v_R3_74_out0;
wire  [15:0] v_R3_75_out0;
wire  [15:0] v_RAM0_1680_out0;
wire  [15:0] v_RAM1_13398_out0;
wire  [15:0] v_RAMDOUT_23_out0;
wire  [15:0] v_RAMDOUT_2414_out0;
wire  [15:0] v_RAMDOUT_2415_out0;
wire  [15:0] v_RAMDOUT_24_out0;
wire  [15:0] v_RAMDOUT_3031_out0;
wire  [15:0] v_RAMDOUT_3032_out0;
wire  [15:0] v_RAM_IN_233_out0;
wire  [15:0] v_RAM_IN_234_out0;
wire  [15:0] v_RAM_OUT0_8764_out0;
wire  [15:0] v_RAM_OUT1_2385_out0;
wire  [15:0] v_RAM_OUT_10335_out0;
wire  [15:0] v_RAM_OUT_10336_out0;
wire  [15:0] v_RAM_OUT_11214_out0;
wire  [15:0] v_RAM_OUT_11215_out0;
wire  [15:0] v_RAM_OUT_1751_out0;
wire  [15:0] v_RAM_OUT_1752_out0;
wire  [15:0] v_RAM_OUT_2104_out0;
wire  [15:0] v_RAM_OUT_2105_out0;
wire  [15:0] v_RAM_OUT_2628_out0;
wire  [15:0] v_RAM_OUT_2629_out0;
wire  [15:0] v_RAM_OUT_3033_out0;
wire  [15:0] v_RAM_OUT_3034_out0;
wire  [15:0] v_RDOUT_2787_out0;
wire  [15:0] v_RDOUT_2788_out0;
wire  [15:0] v_RD_3891_out0;
wire  [15:0] v_RD_3892_out0;
wire  [15:0] v_RD_4839_out0;
wire  [15:0] v_RD_4840_out0;
wire  [15:0] v_RD_501_out0;
wire  [15:0] v_RD_502_out0;
wire  [15:0] v_RD_613_out0;
wire  [15:0] v_RD_614_out0;
wire  [15:0] v_RD_FLOATING_2823_out0;
wire  [15:0] v_RD_FLOATING_2824_out0;
wire  [15:0] v_RD_MULTI_45_out0;
wire  [15:0] v_RD_MULTI_46_out0;
wire  [15:0] v_RD_STATUS_10500_out0;
wire  [15:0] v_REGDIN_11041_out0;
wire  [15:0] v_REGDIN_11042_out0;
wire  [15:0] v_REGISTER_INPUT_13270_out0;
wire  [15:0] v_REGISTER_INPUT_13271_out0;
wire  [15:0] v_REGISTER_INPUT_13621_out0;
wire  [15:0] v_REGISTER_INPUT_13622_out0;
wire  [15:0] v_REGISTER_OUTPUT2_2398_out0;
wire  [15:0] v_REGISTER_OUTPUT_3268_out0;
wire  [15:0] v_REGISTER_OUT_10268_out0;
wire  [15:0] v_REGISTER_OUT_10269_out0;
wire  [15:0] v_REGISTE_IN_4490_out0;
wire  [15:0] v_REGISTE_IN_4491_out0;
wire  [15:0] v_RMN_13437_out0;
wire  [15:0] v_RMN_13438_out0;
wire  [15:0] v_RM_11063_out0;
wire  [15:0] v_RM_11064_out0;
wire  [15:0] v_RM_11065_out0;
wire  [15:0] v_RM_11066_out0;
wire  [15:0] v_RM_11067_out0;
wire  [15:0] v_RM_11068_out0;
wire  [15:0] v_RM_11069_out0;
wire  [15:0] v_RM_11070_out0;
wire  [15:0] v_RM_11071_out0;
wire  [15:0] v_RM_11072_out0;
wire  [15:0] v_RM_11073_out0;
wire  [15:0] v_RM_11074_out0;
wire  [15:0] v_RM_11075_out0;
wire  [15:0] v_RM_11076_out0;
wire  [15:0] v_RM_11077_out0;
wire  [15:0] v_RM_11078_out0;
wire  [15:0] v_RM_11079_out0;
wire  [15:0] v_RM_11080_out0;
wire  [15:0] v_RM_11081_out0;
wire  [15:0] v_RM_11082_out0;
wire  [15:0] v_RM_11083_out0;
wire  [15:0] v_RM_11084_out0;
wire  [15:0] v_RM_11085_out0;
wire  [15:0] v_RM_11086_out0;
wire  [15:0] v_RM_11087_out0;
wire  [15:0] v_RM_11088_out0;
wire  [15:0] v_RM_11089_out0;
wire  [15:0] v_RM_11090_out0;
wire  [15:0] v_RM_11091_out0;
wire  [15:0] v_RM_11092_out0;
wire  [15:0] v_RM_11167_out0;
wire  [15:0] v_RM_11168_out0;
wire  [15:0] v_RM_13508_out0;
wire  [15:0] v_RM_13509_out0;
wire  [15:0] v_RM_13597_out0;
wire  [15:0] v_RM_13598_out0;
wire  [15:0] v_RM_13750_out0;
wire  [15:0] v_RM_13751_out0;
wire  [15:0] v_RM_2432_out0;
wire  [15:0] v_RM_2433_out0;
wire  [15:0] v_RM_2912_out0;
wire  [15:0] v_RM_2913_out0;
wire  [15:0] v_RM_3272_out0;
wire  [15:0] v_RM_3273_out0;
wire  [15:0] v_RM_4537_out0;
wire  [15:0] v_RM_4538_out0;
wire  [15:0] v_RM_8731_out0;
wire  [15:0] v_RM_8732_out0;
wire  [15:0] v_RM_MULTI_210_out0;
wire  [15:0] v_RM_MULTI_211_out0;
wire  [15:0] v_RM_MULTI_648_out0;
wire  [15:0] v_RM_MULTI_649_out0;
wire  [15:0] v_STATUS_REGISTER_10359_out0;
wire  [15:0] v_STATUS_REGISTER_13778_out0;
wire  [15:0] v_STATUS_REGISTER_185_out0;
wire  [15:0] v_STATUS_REGISTER_2866_out0;
wire  [15:0] v_STATUS_REGISTER_2867_out0;
wire  [15:0] v_STATUS_REGISTER_5858_out0;
wire  [15:0] v_STATUS_REGISTER_5859_out0;
wire  [15:0] v_SUM1_13213_out0;
wire  [15:0] v_SUM1_13214_out0;
wire  [15:0] v_XOR1_11246_out0;
wire  [15:0] v_XOR1_11247_out0;
wire  [15:0] v_XOR2_4486_out0;
wire  [15:0] v_XOR2_4487_out0;
wire  [15:0] v_XOR3_13599_out0;
wire  [15:0] v_XOR3_13600_out0;
wire  [15:0] v__10333_out0;
wire  [15:0] v__10334_out0;
wire  [15:0] v__10449_out0;
wire  [15:0] v__10450_out0;
wire  [15:0] v__10504_out0;
wire  [15:0] v__10505_out0;
wire  [15:0] v__10532_out0;
wire  [15:0] v__10814_out0;
wire  [15:0] v__10815_out0;
wire  [15:0] v__10946_out0;
wire  [15:0] v__10947_out0;
wire  [15:0] v__10948_out0;
wire  [15:0] v__10949_out0;
wire  [15:0] v__10950_out0;
wire  [15:0] v__10951_out0;
wire  [15:0] v__10952_out0;
wire  [15:0] v__10953_out0;
wire  [15:0] v__10954_out0;
wire  [15:0] v__10955_out0;
wire  [15:0] v__10956_out0;
wire  [15:0] v__10957_out0;
wire  [15:0] v__10958_out0;
wire  [15:0] v__10959_out0;
wire  [15:0] v__10960_out0;
wire  [15:0] v__10961_out0;
wire  [15:0] v__10962_out0;
wire  [15:0] v__10963_out0;
wire  [15:0] v__10964_out0;
wire  [15:0] v__10965_out0;
wire  [15:0] v__10966_out0;
wire  [15:0] v__10967_out0;
wire  [15:0] v__10968_out0;
wire  [15:0] v__10969_out0;
wire  [15:0] v__10970_out0;
wire  [15:0] v__10971_out0;
wire  [15:0] v__10972_out0;
wire  [15:0] v__10973_out0;
wire  [15:0] v__10974_out0;
wire  [15:0] v__10975_out0;
wire  [15:0] v__11229_out0;
wire  [15:0] v__11230_out0;
wire  [15:0] v__1172_out0;
wire  [15:0] v__1173_out0;
wire  [15:0] v__1209_out0;
wire  [15:0] v__1210_out0;
wire  [15:0] v__1211_out0;
wire  [15:0] v__1212_out0;
wire  [15:0] v__1213_out0;
wire  [15:0] v__1214_out0;
wire  [15:0] v__124_out0;
wire  [15:0] v__125_out0;
wire  [15:0] v__13275_out0;
wire  [15:0] v__13276_out0;
wire  [15:0] v__13482_out0;
wire  [15:0] v__13483_out0;
wire  [15:0] v__167_out0;
wire  [15:0] v__168_out0;
wire  [15:0] v__1867_out0;
wire  [15:0] v__1868_out0;
wire  [15:0] v__1869_out0;
wire  [15:0] v__1870_out0;
wire  [15:0] v__2678_out0;
wire  [15:0] v__2679_out0;
wire  [15:0] v__2791_out0;
wire  [15:0] v__2792_out0;
wire  [15:0] v__3178_out0;
wire  [15:0] v__3179_out0;
wire  [15:0] v__333_out0;
wire  [15:0] v__334_out0;
wire  [15:0] v__403_out0;
wire  [15:0] v__404_out0;
wire  [15:0] v__4660_out0;
wire  [15:0] v__4661_out0;
wire  [15:0] v__4709_out0;
wire  [15:0] v__4710_out0;
wire  [15:0] v__6870_out0;
wire  [15:0] v__6871_out0;
wire  [15:0] v__7081_out0;
wire  [15:0] v__7082_out0;
wire  [15:0] v__7120_out0;
wire  [15:0] v__7121_out0;
wire  [15:0] v__7124_out0;
wire  [15:0] v__7125_out0;
wire  [15:0] v__7179_out0;
wire  [15:0] v__7180_out0;
wire  [15:0] v__7638_out0;
wire  [15:0] v__7639_out0;
wire  [15:0] v__7640_out0;
wire  [15:0] v__7641_out0;
wire  [15:0] v__8697_out0;
wire  [15:0] v__8698_out0;
wire  [15:0] v__9791_out0;
wire  [15:0] v__9792_out0;
wire  [15:0] v_data_ram_1818_out0;
wire  [1:0] v_4BITCOUNTER_317_out0;
wire  [1:0] v_4BITCOUNTER_318_out0;
wire  [1:0] v_4BITCOUNTER_319_out0;
wire  [1:0] v_4BITCOUNTER_320_out0;
wire  [1:0] v_AD1_13774_out0;
wire  [1:0] v_AD1_13775_out0;
wire  [1:0] v_AD2_10699_out0;
wire  [1:0] v_AD2_10700_out0;
wire  [1:0] v_AD3_10482_out0;
wire  [1:0] v_AD3_10483_out0;
wire  [1:0] v_AD3_13272_out0;
wire  [1:0] v_AD3_13273_out0;
wire  [1:0] v_AD3_8671_out0;
wire  [1:0] v_AD3_8672_out0;
wire  [1:0] v_C1_11292_out0;
wire  [1:0] v_C1_11293_out0;
wire  [1:0] v_C1_3205_out0;
wire  [1:0] v_C1_3206_out0;
wire  [1:0] v_C1_6793_out0;
wire  [1:0] v_C1_6794_out0;
wire  [1:0] v_C5_10356_out0;
wire  [1:0] v_D_2108_out0;
wire  [1:0] v_D_2109_out0;
wire  [1:0] v_D_623_out0;
wire  [1:0] v_D_624_out0;
wire  [1:0] v_D_8752_out0;
wire  [1:0] v_D_8753_out0;
wire  [1:0] v_MUX1_11061_out0;
wire  [1:0] v_MUX1_534_out0;
wire  [1:0] v_MUX1_535_out0;
wire  [1:0] v_MUX2_1145_out0;
wire  [1:0] v_MUX2_1146_out0;
wire  [1:0] v_M_4701_out0;
wire  [1:0] v_M_4702_out0;
wire  [1:0] v_M_7177_out0;
wire  [1:0] v_M_7178_out0;
wire  [1:0] v_NOTUSED_2589_out0;
wire  [1:0] v_NOTUSED_2590_out0;
wire  [1:0] v_NOTUSED_445_out0;
wire  [1:0] v_NOTUSED_446_out0;
wire  [1:0] v_NOTUSED_447_out0;
wire  [1:0] v_NOTUSED_448_out0;
wire  [1:0] v_Q_10618_out0;
wire  [1:0] v_Q_1153_out0;
wire  [1:0] v_Q_1154_out0;
wire  [1:0] v_Q_13510_out0;
wire  [1:0] v_RD_10522_out0;
wire  [1:0] v_RD_10523_out0;
wire  [1:0] v_ROR_66_out0;
wire  [1:0] v_ROR_67_out0;
wire  [1:0] v_SHIFT_10615_out0;
wire  [1:0] v_SHIFT_10616_out0;
wire  [1:0] v_SHIFT_8661_out0;
wire  [1:0] v_SHIFT_8662_out0;
wire  [1:0] v_SR_10607_out0;
wire  [1:0] v_SR_10608_out0;
wire  [1:0] v_SR_1956_out0;
wire  [1:0] v_SR_1957_out0;
wire  [1:0] v_SR_371_out0;
wire  [1:0] v_SR_372_out0;
wire  [1:0] v_SR_542_out0;
wire  [1:0] v_SR_543_out0;
wire  [1:0] v_UNUSED_11244_out0;
wire  [1:0] v_UNUSED_11245_out0;
wire  [1:0] v__10287_out0;
wire  [1:0] v__10288_out0;
wire  [1:0] v__10289_out0;
wire  [1:0] v__10290_out0;
wire  [1:0] v__10791_out0;
wire  [1:0] v__10792_out0;
wire  [1:0] v__11049_out1;
wire  [1:0] v__11050_out1;
wire  [1:0] v__11057_out0;
wire  [1:0] v__11058_out0;
wire  [1:0] v__11163_out0;
wire  [1:0] v__11164_out0;
wire  [1:0] v__1140_out0;
wire  [1:0] v__1141_out0;
wire  [1:0] v__13261_out0;
wire  [1:0] v__13262_out0;
wire  [1:0] v__13263_out0;
wire  [1:0] v__13264_out0;
wire  [1:0] v__13550_out0;
wire  [1:0] v__13551_out0;
wire  [1:0] v__13770_out0;
wire  [1:0] v__13771_out0;
wire  [1:0] v__13772_out0;
wire  [1:0] v__13773_out0;
wire  [1:0] v__1707_out0;
wire  [1:0] v__1708_out0;
wire  [1:0] v__1951_out0;
wire  [1:0] v__1952_out0;
wire  [1:0] v__1953_out0;
wire  [1:0] v__1954_out0;
wire  [1:0] v__2599_out0;
wire  [1:0] v__2600_out0;
wire  [1:0] v__2887_out0;
wire  [1:0] v__2888_out0;
wire  [1:0] v__2945_out0;
wire  [1:0] v__2946_out0;
wire  [1:0] v__2947_out0;
wire  [1:0] v__2948_out0;
wire  [1:0] v__3215_out0;
wire  [1:0] v__3216_out0;
wire  [1:0] v__3217_out0;
wire  [1:0] v__3218_out0;
wire  [1:0] v__3223_out0;
wire  [1:0] v__3224_out0;
wire  [1:0] v__3278_out0;
wire  [1:0] v__3279_out0;
wire  [1:0] v__3280_out0;
wire  [1:0] v__3281_out0;
wire  [1:0] v__386_out0;
wire  [1:0] v__387_out0;
wire  [1:0] v__388_out0;
wire  [1:0] v__389_out0;
wire  [1:0] v__399_out0;
wire  [1:0] v__400_out0;
wire  [1:0] v__401_out0;
wire  [1:0] v__402_out0;
wire  [1:0] v__4483_out0;
wire  [1:0] v__4484_out0;
wire  [1:0] v__4547_out0;
wire  [1:0] v__4782_out0;
wire  [1:0] v__4783_out0;
wire  [1:0] v__4784_out0;
wire  [1:0] v__4785_out0;
wire  [1:0] v__4786_out0;
wire  [1:0] v__4787_out0;
wire  [1:0] v__4788_out0;
wire  [1:0] v__4789_out0;
wire  [1:0] v__4790_out0;
wire  [1:0] v__4791_out0;
wire  [1:0] v__4792_out0;
wire  [1:0] v__4793_out0;
wire  [1:0] v__4794_out0;
wire  [1:0] v__4795_out0;
wire  [1:0] v__4796_out0;
wire  [1:0] v__4797_out0;
wire  [1:0] v__4798_out0;
wire  [1:0] v__4799_out0;
wire  [1:0] v__4800_out0;
wire  [1:0] v__4801_out0;
wire  [1:0] v__4802_out0;
wire  [1:0] v__4803_out0;
wire  [1:0] v__4804_out0;
wire  [1:0] v__4805_out0;
wire  [1:0] v__4806_out0;
wire  [1:0] v__4807_out0;
wire  [1:0] v__4808_out0;
wire  [1:0] v__4809_out0;
wire  [1:0] v__4810_out0;
wire  [1:0] v__4811_out0;
wire  [1:0] v__4816_out0;
wire  [1:0] v__4817_out0;
wire  [1:0] v__533_out0;
wire  [1:0] v__627_out0;
wire  [1:0] v__628_out0;
wire  [1:0] v__7135_out0;
wire  [1:0] v__7136_out0;
wire  [1:0] v__7137_out0;
wire  [1:0] v__7138_out0;
wire  [1:0] v__7183_out0;
wire  [1:0] v__7184_out0;
wire  [1:0] v__7185_out0;
wire  [1:0] v__7186_out0;
wire  [2:0] v_C1_2716_out0;
wire  [2:0] v_C2_11233_out0;
wire  [2:0] v_C3_10853_out0;
wire  [2:0] v_C4_1201_out0;
wire  [2:0] v_OP_11223_out0;
wire  [2:0] v_OP_11224_out0;
wire  [2:0] v_OP_621_out0;
wire  [2:0] v_OP_622_out0;
wire  [2:0] v__13253_out0;
wire  [2:0] v__13254_out0;
wire  [2:0] v__1716_out0;
wire  [2:0] v__1717_out0;
wire  [2:0] v__2386_out0;
wire  [2:0] v__2387_out0;
wire  [2:0] v__2552_out0;
wire  [2:0] v__2553_out0;
wire  [2:0] v__2554_out0;
wire  [2:0] v__2555_out0;
wire  [2:0] v__2556_out0;
wire  [2:0] v__2557_out0;
wire  [2:0] v__2558_out0;
wire  [2:0] v__2559_out0;
wire  [2:0] v__2560_out0;
wire  [2:0] v__2561_out0;
wire  [2:0] v__2562_out0;
wire  [2:0] v__2563_out0;
wire  [2:0] v__2564_out0;
wire  [2:0] v__2565_out0;
wire  [2:0] v__2566_out0;
wire  [2:0] v__2567_out0;
wire  [2:0] v__2568_out0;
wire  [2:0] v__2569_out0;
wire  [2:0] v__2570_out0;
wire  [2:0] v__2571_out0;
wire  [2:0] v__2572_out0;
wire  [2:0] v__2573_out0;
wire  [2:0] v__2574_out0;
wire  [2:0] v__2575_out0;
wire  [2:0] v__2576_out0;
wire  [2:0] v__2577_out0;
wire  [2:0] v__2578_out0;
wire  [2:0] v__2579_out0;
wire  [2:0] v__2580_out0;
wire  [2:0] v__2581_out0;
wire  [2:0] v__2680_out1;
wire  [2:0] v__2681_out1;
wire  [2:0] v__2960_out0;
wire  [2:0] v__2961_out0;
wire  [2:0] v__2962_out0;
wire  [2:0] v__2963_out0;
wire  [2:0] v__4_out0;
wire  [2:0] v__5_out0;
wire  [2:0] v__9804_out0;
wire  [2:0] v__9805_out0;
wire  [2:0] v__9806_out0;
wire  [2:0] v__9807_out0;
wire  [31:0] v_32BITPRODUCT_12249_out0;
wire  [31:0] v_32BITPRODUCT_12250_out0;
wire  [31:0] v_32BITPRODUCT_82_out0;
wire  [31:0] v_32BITPRODUCT_83_out0;
wire  [31:0] v_32BIT_MULTI_1183_out0;
wire  [31:0] v_32BIT_MULTI_1184_out0;
wire  [31:0] v_FLOATING_MULTI_7697_out0;
wire  [31:0] v_FLOATING_MULTI_7698_out0;
wire  [31:0] v__212_out0;
wire  [31:0] v__213_out0;
wire  [3:0] v_8BITCOUNTER_13281_out0;
wire  [3:0] v_8BITCOUNTER_13282_out0;
wire  [3:0] v_8BITCOUNTER_13283_out0;
wire  [3:0] v_8BITCOUNTER_13284_out0;
wire  [3:0] v_BIN_5853_out0;
wire  [3:0] v_BIN_5854_out0;
wire  [3:0] v_B_10793_out0;
wire  [3:0] v_B_10794_out0;
wire  [3:0] v_B_1155_out0;
wire  [3:0] v_B_1156_out0;
wire  [3:0] v_B_273_out0;
wire  [3:0] v_B_274_out0;
wire  [3:0] v_C1_10305_out0;
wire  [3:0] v_C1_10306_out0;
wire  [3:0] v_C1_2005_out0;
wire  [3:0] v_C1_2006_out0;
wire  [3:0] v_C1_6919_out0;
wire  [3:0] v_C1_6920_out0;
wire  [3:0] v_MUX1_2409_out0;
wire  [3:0] v_MUX1_2410_out0;
wire  [3:0] v_NOTUSED1_1897_out0;
wire  [3:0] v_NOTUSED1_1898_out0;
wire  [3:0] v_NOTUSED_10540_out0;
wire  [3:0] v_NOTUSED_10541_out0;
wire  [3:0] v_NOTUSED_13265_out0;
wire  [3:0] v_NOTUSED_13266_out0;
wire  [3:0] v_NOTUSED_9800_out0;
wire  [3:0] v_NOTUSED_9801_out0;
wire  [3:0] v_NOTUSE_2399_out0;
wire  [3:0] v_NOTUSE_2400_out0;
wire  [3:0] v_N_7642_out0;
wire  [3:0] v_N_7643_out0;
wire  [3:0] v_RAM_ADD_BYTE0_13382_out0;
wire  [3:0] v_RAM_ADD_BYTE0_13383_out0;
wire  [3:0] v_SEL1_5798_out0;
wire  [3:0] v_SEL1_5799_out0;
wire  [3:0] v_UNUSED_13431_out0;
wire  [3:0] v_UNUSED_13432_out0;
wire  [3:0] v__10372_out0;
wire  [3:0] v__10373_out0;
wire  [3:0] v__10374_out0;
wire  [3:0] v__10375_out0;
wire  [3:0] v__113_out0;
wire  [3:0] v__1140_out1;
wire  [3:0] v__1141_out1;
wire  [3:0] v__114_out0;
wire  [3:0] v__115_out0;
wire  [3:0] v__116_out0;
wire  [3:0] v__13291_out0;
wire  [3:0] v__13292_out0;
wire  [3:0] v__13317_out0;
wire  [3:0] v__13317_out1;
wire  [3:0] v__13318_out0;
wire  [3:0] v__13318_out1;
wire  [3:0] v__13337_out0;
wire  [3:0] v__1673_out0;
wire  [3:0] v__1813_out0;
wire  [3:0] v__2146_out0;
wire  [3:0] v__2147_out0;
wire  [3:0] v__224_out1;
wire  [3:0] v__225_out1;
wire  [3:0] v__2345_out0;
wire  [3:0] v__2346_out0;
wire  [3:0] v__2347_out0;
wire  [3:0] v__2348_out0;
wire  [3:0] v__2411_out1;
wire  [3:0] v__2412_out1;
wire  [3:0] v__2437_out0;
wire  [3:0] v__2438_out0;
wire  [3:0] v__2536_out0;
wire  [3:0] v__2773_out0;
wire  [3:0] v__2774_out0;
wire  [3:0] v__2775_out0;
wire  [3:0] v__2776_out0;
wire  [3:0] v__2968_out0;
wire  [3:0] v__2969_out0;
wire  [3:0] v__3035_out1;
wire  [3:0] v__3036_out1;
wire  [3:0] v__3942_out0;
wire  [3:0] v__3943_out0;
wire  [3:0] v__4488_out0;
wire  [3:0] v__4489_out0;
wire  [3:0] v__449_out0;
wire  [3:0] v__450_out0;
wire  [3:0] v__451_out0;
wire  [3:0] v__4529_out0;
wire  [3:0] v__452_out0;
wire  [3:0] v__4530_out0;
wire  [3:0] v__4585_out0;
wire  [3:0] v__4586_out0;
wire  [3:0] v__4703_out0;
wire  [3:0] v__4704_out0;
wire  [3:0] v__5846_out1;
wire  [3:0] v__5847_out1;
wire  [3:0] v__7032_out0;
wire  [3:0] v__7033_out0;
wire  [3:0] v__7034_out0;
wire  [3:0] v__7035_out0;
wire  [3:0] v__7036_out0;
wire  [3:0] v__7037_out0;
wire  [3:0] v__7038_out0;
wire  [3:0] v__7039_out0;
wire  [3:0] v__7040_out0;
wire  [3:0] v__7041_out0;
wire  [3:0] v__7042_out0;
wire  [3:0] v__7043_out0;
wire  [3:0] v__7044_out0;
wire  [3:0] v__7045_out0;
wire  [3:0] v__7046_out0;
wire  [3:0] v__7047_out0;
wire  [3:0] v__7048_out0;
wire  [3:0] v__7049_out0;
wire  [3:0] v__7050_out0;
wire  [3:0] v__7051_out0;
wire  [3:0] v__7052_out0;
wire  [3:0] v__7053_out0;
wire  [3:0] v__7054_out0;
wire  [3:0] v__7055_out0;
wire  [3:0] v__7056_out0;
wire  [3:0] v__7057_out0;
wire  [3:0] v__7058_out0;
wire  [3:0] v__7059_out0;
wire  [3:0] v__7060_out0;
wire  [3:0] v__7061_out0;
wire  [3:0] v__7116_out1;
wire  [3:0] v__7117_out1;
wire  [3:0] v__8687_out0;
wire  [3:0] v__8688_out0;
wire  [3:0] v__8689_out0;
wire  [3:0] v__8690_out0;
wire  [4:0] v_0B00001_10554_out0;
wire  [4:0] v_0B00001_10555_out0;
wire  [4:0] v_A7_2719_out0;
wire  [4:0] v_A7_2720_out0;
wire  [4:0] v_B_3946_out0;
wire  [4:0] v_B_3947_out0;
wire  [4:0] v_C10_11248_out0;
wire  [4:0] v_C10_11249_out0;
wire  [4:0] v_C14_10795_out0;
wire  [4:0] v_C14_10796_out0;
wire  [4:0] v_C1_10313_out0;
wire  [4:0] v_C1_10314_out0;
wire  [4:0] v_C1_10315_out0;
wire  [4:0] v_C1_10316_out0;
wire  [4:0] v_C4_2593_out0;
wire  [4:0] v_C4_2594_out0;
wire  [4:0] v_C8_2758_out0;
wire  [4:0] v_C8_2759_out0;
wire  [4:0] v_EXP_2441_out0;
wire  [4:0] v_EXP_2442_out0;
wire  [4:0] v_EXP_2907_out0;
wire  [4:0] v_EXP_2908_out0;
wire  [4:0] v_EXP_ANS_10487_out0;
wire  [4:0] v_EXP_ANS_10488_out0;
wire  [4:0] v_EXP_ANS_10860_out0;
wire  [4:0] v_EXP_ANS_10861_out0;
wire  [4:0] v_EXP_ANS_11059_out0;
wire  [4:0] v_EXP_ANS_11060_out0;
wire  [4:0] v_EXP_ANS_13748_out0;
wire  [4:0] v_EXP_ANS_13749_out0;
wire  [4:0] v_EXP_ANS_2008_out0;
wire  [4:0] v_EXP_ANS_2009_out0;
wire  [4:0] v_EXP_PRE_ANS_10765_out0;
wire  [4:0] v_EXP_PRE_ANS_10766_out0;
wire  [4:0] v_EXP_RD_5855_out0;
wire  [4:0] v_EXP_RD_5856_out0;
wire  [4:0] v_EXP_RM_4743_out0;
wire  [4:0] v_EXP_RM_4744_out0;
wire  [4:0] v_K_2636_out0;
wire  [4:0] v_K_2637_out0;
wire  [4:0] v_K_5792_out0;
wire  [4:0] v_K_5793_out0;
wire  [4:0] v_MUX11_86_out0;
wire  [4:0] v_MUX11_87_out0;
wire  [4:0] v_MUX12_13783_out0;
wire  [4:0] v_MUX12_13784_out0;
wire  [4:0] v_MUX13_13647_out0;
wire  [4:0] v_MUX13_13648_out0;
wire  [4:0] v_MUX4_275_out0;
wire  [4:0] v_MUX4_276_out0;
wire  [4:0] v_MUX7_4481_out0;
wire  [4:0] v_MUX7_4482_out0;
wire  [4:0] v_OP2_EXP_10383_out0;
wire  [4:0] v_OP2_EXP_10384_out0;
wire  [4:0] v_OP2_EXP_2548_out0;
wire  [4:0] v_OP2_EXP_2549_out0;
wire  [4:0] v_OP2_EXP_536_out0;
wire  [4:0] v_OP2_EXP_537_out0;
wire  [4:0] v_RD_EXP_2601_out0;
wire  [4:0] v_RD_EXP_2602_out0;
wire  [4:0] v_RD_EXP_3951_out0;
wire  [4:0] v_RD_EXP_3952_out0;
wire  [4:0] v_RD_EXP_8846_out0;
wire  [4:0] v_RD_EXP_8847_out0;
wire  [4:0] v_SEL1_2917_out0;
wire  [4:0] v_SEL1_2918_out0;
wire  [4:0] v_SEL2_13327_out0;
wire  [4:0] v_SEL2_13328_out0;
wire  [4:0] v_SEL3_390_out0;
wire  [4:0] v_SEL3_391_out0;
wire  [4:0] v_SEL4_5790_out0;
wire  [4:0] v_SEL4_5791_out0;
wire  [4:0] v_SHIFT_AMOUNT_226_out0;
wire  [4:0] v_SHIFT_AMOUNT_227_out0;
wire  [4:0] v_SHIFT_AMOUNT_4715_out0;
wire  [4:0] v_SHIFT_AMOUNT_4716_out0;
wire  [4:0] v__13518_out0;
wire  [4:0] v__13519_out0;
wire  [4:0] v__13520_out0;
wire  [4:0] v__13521_out0;
wire  [4:0] v__13522_out0;
wire  [4:0] v__13523_out0;
wire  [4:0] v__13524_out0;
wire  [4:0] v__13525_out0;
wire  [4:0] v__13526_out0;
wire  [4:0] v__13527_out0;
wire  [4:0] v__13528_out0;
wire  [4:0] v__13529_out0;
wire  [4:0] v__13530_out0;
wire  [4:0] v__13531_out0;
wire  [4:0] v__13532_out0;
wire  [4:0] v__13533_out0;
wire  [4:0] v__13534_out0;
wire  [4:0] v__13535_out0;
wire  [4:0] v__13536_out0;
wire  [4:0] v__13537_out0;
wire  [4:0] v__13538_out0;
wire  [4:0] v__13539_out0;
wire  [4:0] v__13540_out0;
wire  [4:0] v__13541_out0;
wire  [4:0] v__13542_out0;
wire  [4:0] v__13543_out0;
wire  [4:0] v__13544_out0;
wire  [4:0] v__13545_out0;
wire  [4:0] v__13546_out0;
wire  [4:0] v__13547_out0;
wire  [4:0] v__2392_out0;
wire  [4:0] v__2393_out0;
wire  [4:0] v__2846_out0;
wire  [4:0] v__2847_out0;
wire  [4:0] v__3251_out0;
wire  [4:0] v__3252_out0;
wire  [4:0] v__3253_out0;
wire  [4:0] v__3254_out0;
wire  [4:0] v__5849_out0;
wire  [4:0] v__5850_out0;
wire  [5:0] v_A4_13603_out0;
wire  [5:0] v_A4_13604_out0;
wire  [5:0] v_A5_2638_out0;
wire  [5:0] v_A5_2639_out0;
wire  [5:0] v_A6_3957_out0;
wire  [5:0] v_A6_3958_out0;
wire  [5:0] v_C11_13765_out0;
wire  [5:0] v_C11_13766_out0;
wire  [5:0] v_C12_2113_out0;
wire  [5:0] v_C12_2114_out0;
wire  [5:0] v_C13_405_out0;
wire  [5:0] v_C13_406_out0;
wire  [5:0] v_C9_11159_out0;
wire  [5:0] v_C9_11160_out0;
wire  [5:0] v_EXP_SUM_5844_out0;
wire  [5:0] v_EXP_SUM_5845_out0;
wire  [5:0] v_MUX10_10395_out0;
wire  [5:0] v_MUX10_10396_out0;
wire  [5:0] v_MUX8_4587_out0;
wire  [5:0] v_MUX8_4588_out0;
wire  [5:0] v_MUX9_13486_out0;
wire  [5:0] v_MUX9_13487_out0;
wire  [5:0] v_NEG1_6921_out0;
wire  [5:0] v_NEG1_6922_out0;
wire  [5:0] v_NOTUSED_2698_out0;
wire  [5:0] v_NOTUSED_2699_out0;
wire  [5:0] v_XOR3_2546_out0;
wire  [5:0] v_XOR3_2547_out0;
wire  [5:0] v_XOR4_6960_out0;
wire  [5:0] v_XOR4_6961_out0;
wire  [5:0] v__10262_out0;
wire  [5:0] v__10263_out0;
wire  [5:0] v__10298_out0;
wire  [5:0] v__10299_out0;
wire  [5:0] v__10300_out0;
wire  [5:0] v__10301_out0;
wire  [5:0] v__10490_out0;
wire  [5:0] v__10491_out0;
wire  [5:0] v__10858_out0;
wire  [5:0] v__10859_out0;
wire  [5:0] v__2610_out0;
wire  [5:0] v__2611_out0;
wire  [5:0] v__3311_out0;
wire  [5:0] v__3312_out0;
wire  [5:0] v__3313_out0;
wire  [5:0] v__3314_out0;
wire  [5:0] v__3315_out0;
wire  [5:0] v__3316_out0;
wire  [5:0] v__3317_out0;
wire  [5:0] v__3318_out0;
wire  [5:0] v__3319_out0;
wire  [5:0] v__3320_out0;
wire  [5:0] v__3321_out0;
wire  [5:0] v__3322_out0;
wire  [5:0] v__3323_out0;
wire  [5:0] v__3324_out0;
wire  [5:0] v__3325_out0;
wire  [5:0] v__3326_out0;
wire  [5:0] v__3327_out0;
wire  [5:0] v__3328_out0;
wire  [5:0] v__3329_out0;
wire  [5:0] v__3330_out0;
wire  [5:0] v__3331_out0;
wire  [5:0] v__3332_out0;
wire  [5:0] v__3333_out0;
wire  [5:0] v__3334_out0;
wire  [5:0] v__3335_out0;
wire  [5:0] v__3336_out0;
wire  [5:0] v__3337_out0;
wire  [5:0] v__3338_out0;
wire  [5:0] v__3339_out0;
wire  [5:0] v__3340_out0;
wire  [5:0] v__3897_out1;
wire  [5:0] v__3898_out1;
wire  [5:0] v__56_out0;
wire  [5:0] v__57_out0;
wire  [5:0] v__96_out0;
wire  [5:0] v__97_out0;
wire  [6:0] v__119_out0;
wire  [6:0] v__120_out0;
wire  [6:0] v__121_out0;
wire  [6:0] v__122_out0;
wire  [6:0] v__2959_out1;
wire  [6:0] v__4703_out1;
wire  [6:0] v__4704_out1;
wire  [6:0] v__681_out0;
wire  [6:0] v__682_out0;
wire  [6:0] v__7062_out0;
wire  [6:0] v__7063_out0;
wire  [6:0] v__7147_out0;
wire  [6:0] v__7148_out0;
wire  [6:0] v__7149_out0;
wire  [6:0] v__7150_out0;
wire  [6:0] v__7151_out0;
wire  [6:0] v__7152_out0;
wire  [6:0] v__7153_out0;
wire  [6:0] v__7154_out0;
wire  [6:0] v__7155_out0;
wire  [6:0] v__7156_out0;
wire  [6:0] v__7157_out0;
wire  [6:0] v__7158_out0;
wire  [6:0] v__7159_out0;
wire  [6:0] v__7160_out0;
wire  [6:0] v__7161_out0;
wire  [6:0] v__7162_out0;
wire  [6:0] v__7163_out0;
wire  [6:0] v__7164_out0;
wire  [6:0] v__7165_out0;
wire  [6:0] v__7166_out0;
wire  [6:0] v__7167_out0;
wire  [6:0] v__7168_out0;
wire  [6:0] v__7169_out0;
wire  [6:0] v__7170_out0;
wire  [6:0] v__7171_out0;
wire  [6:0] v__7172_out0;
wire  [6:0] v__7173_out0;
wire  [6:0] v__7174_out0;
wire  [6:0] v__7175_out0;
wire  [6:0] v__7176_out0;
wire  [6:0] v__72_out0;
wire  [6:0] v__73_out0;
wire  [7:0] v_BYTE_RECEIVED_13441_out0;
wire  [7:0] v_BYTE_RECEIVED_13796_out0;
wire  [7:0] v_BYTE_RECEIVED_2231_out0;
wire  [7:0] v_BYTE_RECEIVED_7101_out0;
wire  [7:0] v_BYTE_RECEIVED_7102_out0;
wire  [7:0] v_BYTE_RECEIVED_8819_out0;
wire  [7:0] v_BYTE_RECEIVED_8820_out0;
wire  [7:0] v_C1_10266_out0;
wire  [7:0] v_C1_10267_out0;
wire  [7:0] v_C1_13277_out0;
wire  [7:0] v_C1_13278_out0;
wire  [7:0] v_C1_13446_out0;
wire  [7:0] v_C1_13447_out0;
wire  [7:0] v_MUX1_13260_out0;
wire  [7:0] v_NOTUSED2_41_out0;
wire  [7:0] v_NOTUSED2_42_out0;
wire  [7:0] v_NOTUSED_10564_out0;
wire  [7:0] v_NOTUSED_10565_out0;
wire  [7:0] v_NOTUSED_683_out0;
wire  [7:0] v_NOTUSED_684_out0;
wire  [7:0] v_NOTUSED_68_out0;
wire  [7:0] v_NOTUSED_69_out0;
wire  [7:0] v_OUT_3037_out0;
wire  [7:0] v_RECEIVERSTREAM_7635_out0;
wire  [7:0] v_RECEIVER_STREAM_564_out0;
wire  [7:0] v_REGISTER_TRANSMIT_DATA_12241_out0;
wire  [7:0] v_TRANSIMISSION_DATA_10818_out0;
wire  [7:0] v_TRANSMISSION_DATA2_7014_out0;
wire  [7:0] v_TRANSMIT_DATA_76_out0;
wire  [7:0] v__10376_out0;
wire  [7:0] v__10868_out0;
wire  [7:0] v__10869_out0;
wire  [7:0] v__11132_out0;
wire  [7:0] v__11132_out1;
wire  [7:0] v__11133_out0;
wire  [7:0] v__11133_out1;
wire  [7:0] v__13790_out0;
wire  [7:0] v__13791_out0;
wire  [7:0] v__13792_out0;
wire  [7:0] v__13793_out0;
wire  [7:0] v__2425_out0;
wire  [7:0] v__2437_out1;
wire  [7:0] v__2438_out1;
wire  [7:0] v__2582_out0;
wire  [7:0] v__2582_out1;
wire  [7:0] v__2583_out0;
wire  [7:0] v__2583_out1;
wire  [7:0] v__2680_out0;
wire  [7:0] v__2681_out0;
wire  [7:0] v__2684_out0;
wire  [7:0] v__2685_out0;
wire  [7:0] v__2686_out0;
wire  [7:0] v__2687_out0;
wire  [7:0] v__3040_out0;
wire  [7:0] v__3125_out0;
wire  [7:0] v__3125_out1;
wire  [7:0] v__3126_out0;
wire  [7:0] v__3126_out1;
wire  [7:0] v__4449_out0;
wire  [7:0] v__4450_out0;
wire  [7:0] v__4451_out0;
wire  [7:0] v__4452_out0;
wire  [7:0] v__4749_out0;
wire  [7:0] v__4750_out0;
wire  [7:0] v__4751_out0;
wire  [7:0] v__4752_out0;
wire  [7:0] v__4753_out0;
wire  [7:0] v__4754_out0;
wire  [7:0] v__4755_out0;
wire  [7:0] v__4756_out0;
wire  [7:0] v__4757_out0;
wire  [7:0] v__4758_out0;
wire  [7:0] v__4759_out0;
wire  [7:0] v__4760_out0;
wire  [7:0] v__4761_out0;
wire  [7:0] v__4762_out0;
wire  [7:0] v__4763_out0;
wire  [7:0] v__4764_out0;
wire  [7:0] v__4765_out0;
wire  [7:0] v__4766_out0;
wire  [7:0] v__4767_out0;
wire  [7:0] v__4768_out0;
wire  [7:0] v__4769_out0;
wire  [7:0] v__4770_out0;
wire  [7:0] v__4771_out0;
wire  [7:0] v__4772_out0;
wire  [7:0] v__4773_out0;
wire  [7:0] v__4774_out0;
wire  [7:0] v__4775_out0;
wire  [7:0] v__4776_out0;
wire  [7:0] v__4777_out0;
wire  [7:0] v__4778_out0;
wire  [7:0] v__636_out0;
wire  [7:0] v__637_out0;
wire  [7:0] v__8673_out0;
wire  [7:0] v__8673_out1;
wire  [7:0] v__8674_out0;
wire  [7:0] v__8674_out1;
wire  [7:0] v__8681_out0;
wire  [7:0] v__8682_out0;
wire  [7:0] v_split_3196_out0;
wire  [7:0] v_split_3196_out1;
wire  [8:0] v_SEL6_3991_out0;
wire  [8:0] v_SEL6_3992_out0;
wire  [8:0] v__13550_out1;
wire  [8:0] v__13551_out1;
wire  [8:0] v__2838_out0;
wire  [8:0] v__2839_out0;
wire  [8:0] v__43_out0;
wire  [8:0] v__44_out0;
wire  [8:0] v__4526_out0;
wire  [8:0] v__4527_out0;
wire  [8:0] v__464_out0;
wire  [8:0] v__465_out0;
wire  [8:0] v__466_out0;
wire  [8:0] v__467_out0;
wire  [8:0] v__6926_out0;
wire  [8:0] v__6927_out0;
wire  [8:0] v__6928_out0;
wire  [8:0] v__6929_out0;
wire  [8:0] v__6930_out0;
wire  [8:0] v__6931_out0;
wire  [8:0] v__6932_out0;
wire  [8:0] v__6933_out0;
wire  [8:0] v__6934_out0;
wire  [8:0] v__6935_out0;
wire  [8:0] v__6936_out0;
wire  [8:0] v__6937_out0;
wire  [8:0] v__6938_out0;
wire  [8:0] v__6939_out0;
wire  [8:0] v__6940_out0;
wire  [8:0] v__6941_out0;
wire  [8:0] v__6942_out0;
wire  [8:0] v__6943_out0;
wire  [8:0] v__6944_out0;
wire  [8:0] v__6945_out0;
wire  [8:0] v__6946_out0;
wire  [8:0] v__6947_out0;
wire  [8:0] v__6948_out0;
wire  [8:0] v__6949_out0;
wire  [8:0] v__6950_out0;
wire  [8:0] v__6951_out0;
wire  [8:0] v__6952_out0;
wire  [8:0] v__6953_out0;
wire  [8:0] v__6954_out0;
wire  [8:0] v__6955_out0;
wire  [8:0] v__7704_out0;
wire  [8:0] v__7705_out0;
wire  [9:0] v_MUX4_10357_out0;
wire  [9:0] v_MUX4_10358_out0;
wire  [9:0] v_MUX6_10350_out0;
wire  [9:0] v_MUX6_10351_out0;
wire  [9:0] v_OP2_SIG_13301_out0;
wire  [9:0] v_OP2_SIG_13302_out0;
wire  [9:0] v_RD_SIG_1769_out0;
wire  [9:0] v_RD_SIG_1770_out0;
wire  [9:0] v_SEL4_11225_out0;
wire  [9:0] v_SEL4_11226_out0;
wire  [9:0] v_SEL5_8767_out0;
wire  [9:0] v_SEL5_8768_out0;
wire  [9:0] v_SEL6_103_out0;
wire  [9:0] v_SEL6_104_out0;
wire  [9:0] v_SEL9_13753_out0;
wire  [9:0] v_SEL9_13754_out0;
wire  [9:0] v_SIG_ANS_10296_out0;
wire  [9:0] v_SIG_ANS_10297_out0;
wire  [9:0] v_SIG_ANS_2335_out0;
wire  [9:0] v_SIG_ANS_2336_out0;
wire  [9:0] v_SIG_ANS_3276_out0;
wire  [9:0] v_SIG_ANS_3277_out0;
wire  [9:0] v_SIG_ANS_439_out0;
wire  [9:0] v_SIG_ANS_440_out0;
wire  [9:0] v_SIG_RD_11298_out0;
wire  [9:0] v_SIG_RD_11299_out0;
wire  [9:0] v_SIG_RM_1767_out0;
wire  [9:0] v_SIG_RM_1768_out0;
wire  [9:0] v__10775_out0;
wire  [9:0] v__10776_out0;
wire  [9:0] v__10806_out0;
wire  [9:0] v__10807_out0;
wire  [9:0] v__2649_out0;
wire  [9:0] v__2650_out0;
wire  [9:0] v__3897_out0;
wire  [9:0] v__3898_out0;
wire  [9:0] v__3907_out1;
wire  [9:0] v__3908_out1;
wire  [9:0] v__422_out0;
wire  [9:0] v__423_out0;
wire  [9:0] v__424_out0;
wire  [9:0] v__425_out0;
wire  [9:0] v__5802_out0;
wire  [9:0] v__5803_out0;
wire  [9:0] v__5804_out0;
wire  [9:0] v__5805_out0;
wire  [9:0] v__5806_out0;
wire  [9:0] v__5807_out0;
wire  [9:0] v__5808_out0;
wire  [9:0] v__5809_out0;
wire  [9:0] v__5810_out0;
wire  [9:0] v__5811_out0;
wire  [9:0] v__5812_out0;
wire  [9:0] v__5813_out0;
wire  [9:0] v__5814_out0;
wire  [9:0] v__5815_out0;
wire  [9:0] v__5816_out0;
wire  [9:0] v__5817_out0;
wire  [9:0] v__5818_out0;
wire  [9:0] v__5819_out0;
wire  [9:0] v__5820_out0;
wire  [9:0] v__5821_out0;
wire  [9:0] v__5822_out0;
wire  [9:0] v__5823_out0;
wire  [9:0] v__5824_out0;
wire  [9:0] v__5825_out0;
wire  [9:0] v__5826_out0;
wire  [9:0] v__5827_out0;
wire  [9:0] v__5828_out0;
wire  [9:0] v__5829_out0;
wire  [9:0] v__5830_out0;
wire  [9:0] v__5831_out0;
wire  [9:0] v__8677_out0;
wire  [9:0] v__8678_out0;
wire v_0_10706_out0;
wire v_0_10707_out0;
wire v_0_3022_out0;
wire v_0_3023_out0;
wire v_1_3817_out0;
wire v_1_3818_out0;
wire v_2_1763_out0;
wire v_2_1764_out0;
wire v_2_7072_out0;
wire v_3_13619_out0;
wire v_3_13620_out0;
wire v_9_13623_out0;
wire v_9_13624_out0;
wire v_9_13625_out0;
wire v_9_13626_out0;
wire v_9_1700_out0;
wire v_9_1701_out0;
wire v_9_1702_out0;
wire v_9_1703_out0;
wire v_9_417_out0;
wire v_A1_11043_out1;
wire v_A1_3174_out1;
wire v_A1_3175_out1;
wire v_A1_3855_out1;
wire v_A1_3856_out1;
wire v_A1_7019_out1;
wire v_A1_7020_out1;
wire v_A4_11227_out1;
wire v_A4_11228_out1;
wire v_A4_13603_out1;
wire v_A4_13604_out1;
wire v_A5_1901_out1;
wire v_A5_1902_out1;
wire v_A5_2638_out1;
wire v_A5_2639_out1;
wire v_A6_10463_out1;
wire v_A6_10464_out1;
wire v_A6_3957_out1;
wire v_A6_3958_out1;
wire v_A7_2719_out1;
wire v_A7_2720_out1;
wire v_A8_11155_out1;
wire v_A8_11156_out1;
wire v_ADC_10393_out0;
wire v_ADC_10394_out0;
wire v_ADC_13614_out0;
wire v_ADC_13615_out0;
wire v_ADC_1821_out0;
wire v_ADC_1822_out0;
wire v_ADD_11193_out0;
wire v_ADD_11194_out0;
wire v_ADD_4455_out0;
wire v_ADD_4456_out0;
wire v_AND_13556_out0;
wire v_AND_13557_out0;
wire v_AND_3858_out0;
wire v_AND_3859_out0;
wire v_ASR_10366_out0;
wire v_ASR_10367_out0;
wire v_ASR_10566_out0;
wire v_ASR_10567_out0;
wire v_ASR_13713_out0;
wire v_ASR_13714_out0;
wire v_ASR_8754_out0;
wire v_ASR_8755_out0;
wire v_BIT10_7009_out0;
wire v_BIT10_7010_out0;
wire v_BIT_2328_out0;
wire v_BIT_383_out0;
wire v_BIT_6918_out0;
wire v_BIT_IN1_3209_out0;
wire v_BIT_OUT_10705_out0;
wire v_BIT_OUT_13326_out0;
wire v_BIT_OUT_2015_out0;
wire v_BIT_STREAM_IN_13_out0;
wire v_BYTE1_comp1_2443_out0;
wire v_BYTE1_comp1_2444_out0;
wire v_BYTE2_COMP8_7695_out0;
wire v_BYTE2_COMP8_7696_out0;
wire v_BYTERECEIVED_11197_out0;
wire v_BYTE_COMP1_3262_out0;
wire v_BYTE_COMP1_3263_out0;
wire v_BYTE_COMP1_9796_out0;
wire v_BYTE_COMP1_9797_out0;
wire v_BYTE_COMP_10_13611_out0;
wire v_BYTE_COMP_11_1163_out0;
wire v_BYTE_COMP_1_8743_out0;
wire v_BYTE_READY_10558_out0;
wire v_BYTE_READY_10559_out0;
wire v_BYTE_READY_11172_out0;
wire v_BYTE_READY_11173_out0;
wire v_BYTE_READY_13255_out0;
wire v_BYTE_READY_2852_out0;
wire v_BYTE_READY_2853_out0;
wire v_BYTE_READY_7021_out0;
wire v_BYTE_READY_7022_out0;
wire v_C10_1819_out0;
wire v_C10_1820_out0;
wire v_C12_1151_out0;
wire v_C12_1152_out0;
wire v_C14_1674_out0;
wire v_C14_1675_out0;
wire v_C1_10259_out0;
wire v_C1_10789_out0;
wire v_C1_10790_out0;
wire v_C1_436_out0;
wire v_C1_604_out0;
wire v_C1_605_out0;
wire v_C1_8815_out0;
wire v_C1_8816_out0;
wire v_C3_2764_out0;
wire v_C3_4741_out0;
wire v_C3_4742_out0;
wire v_C4_10619_out0;
wire v_C4_90_out0;
wire v_C5_11031_out0;
wire v_C5_13267_out0;
wire v_C6_10317_out0;
wire v_C6_10318_out0;
wire v_C6_1732_out0;
wire v_C7_2271_out0;
wire v_C7_2272_out0;
wire v_C7_3222_out0;
wire v_C9_3029_out0;
wire v_C9_3030_out0;
wire v_CARRY_4862_out0;
wire v_CARRY_4863_out0;
wire v_CARRY_4864_out0;
wire v_CARRY_4865_out0;
wire v_CARRY_4866_out0;
wire v_CARRY_4867_out0;
wire v_CARRY_4868_out0;
wire v_CARRY_4869_out0;
wire v_CARRY_4870_out0;
wire v_CARRY_4871_out0;
wire v_CARRY_4872_out0;
wire v_CARRY_4873_out0;
wire v_CARRY_4874_out0;
wire v_CARRY_4875_out0;
wire v_CARRY_4876_out0;
wire v_CARRY_4877_out0;
wire v_CARRY_4878_out0;
wire v_CARRY_4879_out0;
wire v_CARRY_4880_out0;
wire v_CARRY_4881_out0;
wire v_CARRY_4882_out0;
wire v_CARRY_4883_out0;
wire v_CARRY_4884_out0;
wire v_CARRY_4885_out0;
wire v_CARRY_4886_out0;
wire v_CARRY_4887_out0;
wire v_CARRY_4888_out0;
wire v_CARRY_4889_out0;
wire v_CARRY_4890_out0;
wire v_CARRY_4891_out0;
wire v_CARRY_4892_out0;
wire v_CARRY_4893_out0;
wire v_CARRY_4894_out0;
wire v_CARRY_4895_out0;
wire v_CARRY_4896_out0;
wire v_CARRY_4897_out0;
wire v_CARRY_4898_out0;
wire v_CARRY_4899_out0;
wire v_CARRY_4900_out0;
wire v_CARRY_4901_out0;
wire v_CARRY_4902_out0;
wire v_CARRY_4903_out0;
wire v_CARRY_4904_out0;
wire v_CARRY_4905_out0;
wire v_CARRY_4906_out0;
wire v_CARRY_4907_out0;
wire v_CARRY_4908_out0;
wire v_CARRY_4909_out0;
wire v_CARRY_4910_out0;
wire v_CARRY_4911_out0;
wire v_CARRY_4912_out0;
wire v_CARRY_4913_out0;
wire v_CARRY_4914_out0;
wire v_CARRY_4915_out0;
wire v_CARRY_4916_out0;
wire v_CARRY_4917_out0;
wire v_CARRY_4918_out0;
wire v_CARRY_4919_out0;
wire v_CARRY_4920_out0;
wire v_CARRY_4921_out0;
wire v_CARRY_4922_out0;
wire v_CARRY_4923_out0;
wire v_CARRY_4924_out0;
wire v_CARRY_4925_out0;
wire v_CARRY_4926_out0;
wire v_CARRY_4927_out0;
wire v_CARRY_4928_out0;
wire v_CARRY_4929_out0;
wire v_CARRY_4930_out0;
wire v_CARRY_4931_out0;
wire v_CARRY_4932_out0;
wire v_CARRY_4933_out0;
wire v_CARRY_4934_out0;
wire v_CARRY_4935_out0;
wire v_CARRY_4936_out0;
wire v_CARRY_4937_out0;
wire v_CARRY_4938_out0;
wire v_CARRY_4939_out0;
wire v_CARRY_4940_out0;
wire v_CARRY_4941_out0;
wire v_CARRY_4942_out0;
wire v_CARRY_4943_out0;
wire v_CARRY_4944_out0;
wire v_CARRY_4945_out0;
wire v_CARRY_4946_out0;
wire v_CARRY_4947_out0;
wire v_CARRY_4948_out0;
wire v_CARRY_4949_out0;
wire v_CARRY_4950_out0;
wire v_CARRY_4951_out0;
wire v_CARRY_4952_out0;
wire v_CARRY_4953_out0;
wire v_CARRY_4954_out0;
wire v_CARRY_4955_out0;
wire v_CARRY_4956_out0;
wire v_CARRY_4957_out0;
wire v_CARRY_4958_out0;
wire v_CARRY_4959_out0;
wire v_CARRY_4960_out0;
wire v_CARRY_4961_out0;
wire v_CARRY_4962_out0;
wire v_CARRY_4963_out0;
wire v_CARRY_4964_out0;
wire v_CARRY_4965_out0;
wire v_CARRY_4966_out0;
wire v_CARRY_4967_out0;
wire v_CARRY_4968_out0;
wire v_CARRY_4969_out0;
wire v_CARRY_4970_out0;
wire v_CARRY_4971_out0;
wire v_CARRY_4972_out0;
wire v_CARRY_4973_out0;
wire v_CARRY_4974_out0;
wire v_CARRY_4975_out0;
wire v_CARRY_4976_out0;
wire v_CARRY_4977_out0;
wire v_CARRY_4978_out0;
wire v_CARRY_4979_out0;
wire v_CARRY_4980_out0;
wire v_CARRY_4981_out0;
wire v_CARRY_4982_out0;
wire v_CARRY_4983_out0;
wire v_CARRY_4984_out0;
wire v_CARRY_4985_out0;
wire v_CARRY_4986_out0;
wire v_CARRY_4987_out0;
wire v_CARRY_4988_out0;
wire v_CARRY_4989_out0;
wire v_CARRY_4990_out0;
wire v_CARRY_4991_out0;
wire v_CARRY_4992_out0;
wire v_CARRY_4993_out0;
wire v_CARRY_4994_out0;
wire v_CARRY_4995_out0;
wire v_CARRY_4996_out0;
wire v_CARRY_4997_out0;
wire v_CARRY_4998_out0;
wire v_CARRY_4999_out0;
wire v_CARRY_5000_out0;
wire v_CARRY_5001_out0;
wire v_CARRY_5002_out0;
wire v_CARRY_5003_out0;
wire v_CARRY_5004_out0;
wire v_CARRY_5005_out0;
wire v_CARRY_5006_out0;
wire v_CARRY_5007_out0;
wire v_CARRY_5008_out0;
wire v_CARRY_5009_out0;
wire v_CARRY_5010_out0;
wire v_CARRY_5011_out0;
wire v_CARRY_5012_out0;
wire v_CARRY_5013_out0;
wire v_CARRY_5014_out0;
wire v_CARRY_5015_out0;
wire v_CARRY_5016_out0;
wire v_CARRY_5017_out0;
wire v_CARRY_5018_out0;
wire v_CARRY_5019_out0;
wire v_CARRY_5020_out0;
wire v_CARRY_5021_out0;
wire v_CARRY_5022_out0;
wire v_CARRY_5023_out0;
wire v_CARRY_5024_out0;
wire v_CARRY_5025_out0;
wire v_CARRY_5026_out0;
wire v_CARRY_5027_out0;
wire v_CARRY_5028_out0;
wire v_CARRY_5029_out0;
wire v_CARRY_5030_out0;
wire v_CARRY_5031_out0;
wire v_CARRY_5032_out0;
wire v_CARRY_5033_out0;
wire v_CARRY_5034_out0;
wire v_CARRY_5035_out0;
wire v_CARRY_5036_out0;
wire v_CARRY_5037_out0;
wire v_CARRY_5038_out0;
wire v_CARRY_5039_out0;
wire v_CARRY_5040_out0;
wire v_CARRY_5041_out0;
wire v_CARRY_5042_out0;
wire v_CARRY_5043_out0;
wire v_CARRY_5044_out0;
wire v_CARRY_5045_out0;
wire v_CARRY_5046_out0;
wire v_CARRY_5047_out0;
wire v_CARRY_5048_out0;
wire v_CARRY_5049_out0;
wire v_CARRY_5050_out0;
wire v_CARRY_5051_out0;
wire v_CARRY_5052_out0;
wire v_CARRY_5053_out0;
wire v_CARRY_5054_out0;
wire v_CARRY_5055_out0;
wire v_CARRY_5056_out0;
wire v_CARRY_5057_out0;
wire v_CARRY_5058_out0;
wire v_CARRY_5059_out0;
wire v_CARRY_5060_out0;
wire v_CARRY_5061_out0;
wire v_CARRY_5062_out0;
wire v_CARRY_5063_out0;
wire v_CARRY_5064_out0;
wire v_CARRY_5065_out0;
wire v_CARRY_5066_out0;
wire v_CARRY_5067_out0;
wire v_CARRY_5068_out0;
wire v_CARRY_5069_out0;
wire v_CARRY_5070_out0;
wire v_CARRY_5071_out0;
wire v_CARRY_5072_out0;
wire v_CARRY_5073_out0;
wire v_CARRY_5074_out0;
wire v_CARRY_5075_out0;
wire v_CARRY_5076_out0;
wire v_CARRY_5077_out0;
wire v_CARRY_5078_out0;
wire v_CARRY_5079_out0;
wire v_CARRY_5080_out0;
wire v_CARRY_5081_out0;
wire v_CARRY_5082_out0;
wire v_CARRY_5083_out0;
wire v_CARRY_5084_out0;
wire v_CARRY_5085_out0;
wire v_CARRY_5086_out0;
wire v_CARRY_5087_out0;
wire v_CARRY_5088_out0;
wire v_CARRY_5089_out0;
wire v_CARRY_5090_out0;
wire v_CARRY_5091_out0;
wire v_CARRY_5092_out0;
wire v_CARRY_5093_out0;
wire v_CARRY_5094_out0;
wire v_CARRY_5095_out0;
wire v_CARRY_5096_out0;
wire v_CARRY_5097_out0;
wire v_CARRY_5098_out0;
wire v_CARRY_5099_out0;
wire v_CARRY_5100_out0;
wire v_CARRY_5101_out0;
wire v_CARRY_5102_out0;
wire v_CARRY_5103_out0;
wire v_CARRY_5104_out0;
wire v_CARRY_5105_out0;
wire v_CARRY_5106_out0;
wire v_CARRY_5107_out0;
wire v_CARRY_5108_out0;
wire v_CARRY_5109_out0;
wire v_CARRY_5110_out0;
wire v_CARRY_5111_out0;
wire v_CARRY_5112_out0;
wire v_CARRY_5113_out0;
wire v_CARRY_5114_out0;
wire v_CARRY_5115_out0;
wire v_CARRY_5116_out0;
wire v_CARRY_5117_out0;
wire v_CARRY_5118_out0;
wire v_CARRY_5119_out0;
wire v_CARRY_5120_out0;
wire v_CARRY_5121_out0;
wire v_CARRY_5122_out0;
wire v_CARRY_5123_out0;
wire v_CARRY_5124_out0;
wire v_CARRY_5125_out0;
wire v_CARRY_5126_out0;
wire v_CARRY_5127_out0;
wire v_CARRY_5128_out0;
wire v_CARRY_5129_out0;
wire v_CARRY_5130_out0;
wire v_CARRY_5131_out0;
wire v_CARRY_5132_out0;
wire v_CARRY_5133_out0;
wire v_CARRY_5134_out0;
wire v_CARRY_5135_out0;
wire v_CARRY_5136_out0;
wire v_CARRY_5137_out0;
wire v_CARRY_5138_out0;
wire v_CARRY_5139_out0;
wire v_CARRY_5140_out0;
wire v_CARRY_5141_out0;
wire v_CARRY_5142_out0;
wire v_CARRY_5143_out0;
wire v_CARRY_5144_out0;
wire v_CARRY_5145_out0;
wire v_CARRY_5146_out0;
wire v_CARRY_5147_out0;
wire v_CARRY_5148_out0;
wire v_CARRY_5149_out0;
wire v_CARRY_5150_out0;
wire v_CARRY_5151_out0;
wire v_CARRY_5152_out0;
wire v_CARRY_5153_out0;
wire v_CARRY_5154_out0;
wire v_CARRY_5155_out0;
wire v_CARRY_5156_out0;
wire v_CARRY_5157_out0;
wire v_CARRY_5158_out0;
wire v_CARRY_5159_out0;
wire v_CARRY_5160_out0;
wire v_CARRY_5161_out0;
wire v_CARRY_5162_out0;
wire v_CARRY_5163_out0;
wire v_CARRY_5164_out0;
wire v_CARRY_5165_out0;
wire v_CARRY_5166_out0;
wire v_CARRY_5167_out0;
wire v_CARRY_5168_out0;
wire v_CARRY_5169_out0;
wire v_CARRY_5170_out0;
wire v_CARRY_5171_out0;
wire v_CARRY_5172_out0;
wire v_CARRY_5173_out0;
wire v_CARRY_5174_out0;
wire v_CARRY_5175_out0;
wire v_CARRY_5176_out0;
wire v_CARRY_5177_out0;
wire v_CARRY_5178_out0;
wire v_CARRY_5179_out0;
wire v_CARRY_5180_out0;
wire v_CARRY_5181_out0;
wire v_CARRY_5182_out0;
wire v_CARRY_5183_out0;
wire v_CARRY_5184_out0;
wire v_CARRY_5185_out0;
wire v_CARRY_5186_out0;
wire v_CARRY_5187_out0;
wire v_CARRY_5188_out0;
wire v_CARRY_5189_out0;
wire v_CARRY_5190_out0;
wire v_CARRY_5191_out0;
wire v_CARRY_5192_out0;
wire v_CARRY_5193_out0;
wire v_CARRY_5194_out0;
wire v_CARRY_5195_out0;
wire v_CARRY_5196_out0;
wire v_CARRY_5197_out0;
wire v_CARRY_5198_out0;
wire v_CARRY_5199_out0;
wire v_CARRY_5200_out0;
wire v_CARRY_5201_out0;
wire v_CARRY_5202_out0;
wire v_CARRY_5203_out0;
wire v_CARRY_5204_out0;
wire v_CARRY_5205_out0;
wire v_CARRY_5206_out0;
wire v_CARRY_5207_out0;
wire v_CARRY_5208_out0;
wire v_CARRY_5209_out0;
wire v_CARRY_5210_out0;
wire v_CARRY_5211_out0;
wire v_CARRY_5212_out0;
wire v_CARRY_5213_out0;
wire v_CARRY_5214_out0;
wire v_CARRY_5215_out0;
wire v_CARRY_5216_out0;
wire v_CARRY_5217_out0;
wire v_CARRY_5218_out0;
wire v_CARRY_5219_out0;
wire v_CARRY_5220_out0;
wire v_CARRY_5221_out0;
wire v_CARRY_5222_out0;
wire v_CARRY_5223_out0;
wire v_CARRY_5224_out0;
wire v_CARRY_5225_out0;
wire v_CARRY_5226_out0;
wire v_CARRY_5227_out0;
wire v_CARRY_5228_out0;
wire v_CARRY_5229_out0;
wire v_CARRY_5230_out0;
wire v_CARRY_5231_out0;
wire v_CARRY_5232_out0;
wire v_CARRY_5233_out0;
wire v_CARRY_5234_out0;
wire v_CARRY_5235_out0;
wire v_CARRY_5236_out0;
wire v_CARRY_5237_out0;
wire v_CARRY_5238_out0;
wire v_CARRY_5239_out0;
wire v_CARRY_5240_out0;
wire v_CARRY_5241_out0;
wire v_CARRY_5242_out0;
wire v_CARRY_5243_out0;
wire v_CARRY_5244_out0;
wire v_CARRY_5245_out0;
wire v_CARRY_5246_out0;
wire v_CARRY_5247_out0;
wire v_CARRY_5248_out0;
wire v_CARRY_5249_out0;
wire v_CARRY_5250_out0;
wire v_CARRY_5251_out0;
wire v_CARRY_5252_out0;
wire v_CARRY_5253_out0;
wire v_CARRY_5254_out0;
wire v_CARRY_5255_out0;
wire v_CARRY_5256_out0;
wire v_CARRY_5257_out0;
wire v_CARRY_5258_out0;
wire v_CARRY_5259_out0;
wire v_CARRY_5260_out0;
wire v_CARRY_5261_out0;
wire v_CARRY_5262_out0;
wire v_CARRY_5263_out0;
wire v_CARRY_5264_out0;
wire v_CARRY_5265_out0;
wire v_CARRY_5266_out0;
wire v_CARRY_5267_out0;
wire v_CARRY_5268_out0;
wire v_CARRY_5269_out0;
wire v_CARRY_5270_out0;
wire v_CARRY_5271_out0;
wire v_CARRY_5272_out0;
wire v_CARRY_5273_out0;
wire v_CARRY_5274_out0;
wire v_CARRY_5275_out0;
wire v_CARRY_5276_out0;
wire v_CARRY_5277_out0;
wire v_CARRY_5278_out0;
wire v_CARRY_5279_out0;
wire v_CARRY_5280_out0;
wire v_CARRY_5281_out0;
wire v_CARRY_5282_out0;
wire v_CARRY_5283_out0;
wire v_CARRY_5284_out0;
wire v_CARRY_5285_out0;
wire v_CARRY_5286_out0;
wire v_CARRY_5287_out0;
wire v_CARRY_5288_out0;
wire v_CARRY_5289_out0;
wire v_CARRY_5290_out0;
wire v_CARRY_5291_out0;
wire v_CARRY_5292_out0;
wire v_CARRY_5293_out0;
wire v_CARRY_5294_out0;
wire v_CARRY_5295_out0;
wire v_CARRY_5296_out0;
wire v_CARRY_5297_out0;
wire v_CARRY_5298_out0;
wire v_CARRY_5299_out0;
wire v_CARRY_5300_out0;
wire v_CARRY_5301_out0;
wire v_CARRY_5302_out0;
wire v_CARRY_5303_out0;
wire v_CARRY_5304_out0;
wire v_CARRY_5305_out0;
wire v_CARRY_5306_out0;
wire v_CARRY_5307_out0;
wire v_CARRY_5308_out0;
wire v_CARRY_5309_out0;
wire v_CARRY_5310_out0;
wire v_CARRY_5311_out0;
wire v_CARRY_5312_out0;
wire v_CARRY_5313_out0;
wire v_CARRY_5314_out0;
wire v_CARRY_5315_out0;
wire v_CARRY_5316_out0;
wire v_CARRY_5317_out0;
wire v_CARRY_5318_out0;
wire v_CARRY_5319_out0;
wire v_CARRY_5320_out0;
wire v_CARRY_5321_out0;
wire v_CARRY_5322_out0;
wire v_CARRY_5323_out0;
wire v_CARRY_5324_out0;
wire v_CARRY_5325_out0;
wire v_CARRY_5326_out0;
wire v_CARRY_5327_out0;
wire v_CARRY_5328_out0;
wire v_CARRY_5329_out0;
wire v_CARRY_5330_out0;
wire v_CARRY_5331_out0;
wire v_CARRY_5332_out0;
wire v_CARRY_5333_out0;
wire v_CARRY_5334_out0;
wire v_CARRY_5335_out0;
wire v_CARRY_5336_out0;
wire v_CARRY_5337_out0;
wire v_CARRY_5338_out0;
wire v_CARRY_5339_out0;
wire v_CARRY_5340_out0;
wire v_CARRY_5341_out0;
wire v_CARRY_5342_out0;
wire v_CARRY_5343_out0;
wire v_CARRY_5344_out0;
wire v_CARRY_5345_out0;
wire v_CARRY_5346_out0;
wire v_CARRY_5347_out0;
wire v_CARRY_5348_out0;
wire v_CARRY_5349_out0;
wire v_CARRY_5350_out0;
wire v_CARRY_5351_out0;
wire v_CARRY_5352_out0;
wire v_CARRY_5353_out0;
wire v_CARRY_5354_out0;
wire v_CARRY_5355_out0;
wire v_CARRY_5356_out0;
wire v_CARRY_5357_out0;
wire v_CARRY_5358_out0;
wire v_CARRY_5359_out0;
wire v_CARRY_5360_out0;
wire v_CARRY_5361_out0;
wire v_CARRY_5362_out0;
wire v_CARRY_5363_out0;
wire v_CARRY_5364_out0;
wire v_CARRY_5365_out0;
wire v_CARRY_5366_out0;
wire v_CARRY_5367_out0;
wire v_CARRY_5368_out0;
wire v_CARRY_5369_out0;
wire v_CARRY_5370_out0;
wire v_CARRY_5371_out0;
wire v_CARRY_5372_out0;
wire v_CARRY_5373_out0;
wire v_CARRY_5374_out0;
wire v_CARRY_5375_out0;
wire v_CARRY_5376_out0;
wire v_CARRY_5377_out0;
wire v_CARRY_5378_out0;
wire v_CARRY_5379_out0;
wire v_CARRY_5380_out0;
wire v_CARRY_5381_out0;
wire v_CARRY_5382_out0;
wire v_CARRY_5383_out0;
wire v_CARRY_5384_out0;
wire v_CARRY_5385_out0;
wire v_CARRY_5386_out0;
wire v_CARRY_5387_out0;
wire v_CARRY_5388_out0;
wire v_CARRY_5389_out0;
wire v_CARRY_5390_out0;
wire v_CARRY_5391_out0;
wire v_CARRY_5392_out0;
wire v_CARRY_5393_out0;
wire v_CARRY_5394_out0;
wire v_CARRY_5395_out0;
wire v_CARRY_5396_out0;
wire v_CARRY_5397_out0;
wire v_CARRY_5398_out0;
wire v_CARRY_5399_out0;
wire v_CARRY_5400_out0;
wire v_CARRY_5401_out0;
wire v_CARRY_5402_out0;
wire v_CARRY_5403_out0;
wire v_CARRY_5404_out0;
wire v_CARRY_5405_out0;
wire v_CARRY_5406_out0;
wire v_CARRY_5407_out0;
wire v_CARRY_5408_out0;
wire v_CARRY_5409_out0;
wire v_CARRY_5410_out0;
wire v_CARRY_5411_out0;
wire v_CARRY_5412_out0;
wire v_CARRY_5413_out0;
wire v_CARRY_5414_out0;
wire v_CARRY_5415_out0;
wire v_CARRY_5416_out0;
wire v_CARRY_5417_out0;
wire v_CARRY_5418_out0;
wire v_CARRY_5419_out0;
wire v_CARRY_5420_out0;
wire v_CARRY_5421_out0;
wire v_CARRY_5422_out0;
wire v_CARRY_5423_out0;
wire v_CARRY_5424_out0;
wire v_CARRY_5425_out0;
wire v_CARRY_5426_out0;
wire v_CARRY_5427_out0;
wire v_CARRY_5428_out0;
wire v_CARRY_5429_out0;
wire v_CARRY_5430_out0;
wire v_CARRY_5431_out0;
wire v_CARRY_5432_out0;
wire v_CARRY_5433_out0;
wire v_CARRY_5434_out0;
wire v_CARRY_5435_out0;
wire v_CARRY_5436_out0;
wire v_CARRY_5437_out0;
wire v_CARRY_5438_out0;
wire v_CARRY_5439_out0;
wire v_CARRY_5440_out0;
wire v_CARRY_5441_out0;
wire v_CARRY_5442_out0;
wire v_CARRY_5443_out0;
wire v_CARRY_5444_out0;
wire v_CARRY_5445_out0;
wire v_CARRY_5446_out0;
wire v_CARRY_5447_out0;
wire v_CARRY_5448_out0;
wire v_CARRY_5449_out0;
wire v_CARRY_5450_out0;
wire v_CARRY_5451_out0;
wire v_CARRY_5452_out0;
wire v_CARRY_5453_out0;
wire v_CARRY_5454_out0;
wire v_CARRY_5455_out0;
wire v_CARRY_5456_out0;
wire v_CARRY_5457_out0;
wire v_CARRY_5458_out0;
wire v_CARRY_5459_out0;
wire v_CARRY_5460_out0;
wire v_CARRY_5461_out0;
wire v_CARRY_5462_out0;
wire v_CARRY_5463_out0;
wire v_CARRY_5464_out0;
wire v_CARRY_5465_out0;
wire v_CARRY_5466_out0;
wire v_CARRY_5467_out0;
wire v_CARRY_5468_out0;
wire v_CARRY_5469_out0;
wire v_CARRY_5470_out0;
wire v_CARRY_5471_out0;
wire v_CARRY_5472_out0;
wire v_CARRY_5473_out0;
wire v_CARRY_5474_out0;
wire v_CARRY_5475_out0;
wire v_CARRY_5476_out0;
wire v_CARRY_5477_out0;
wire v_CARRY_5478_out0;
wire v_CARRY_5479_out0;
wire v_CARRY_5480_out0;
wire v_CARRY_5481_out0;
wire v_CARRY_5482_out0;
wire v_CARRY_5483_out0;
wire v_CARRY_5484_out0;
wire v_CARRY_5485_out0;
wire v_CARRY_5486_out0;
wire v_CARRY_5487_out0;
wire v_CARRY_5488_out0;
wire v_CARRY_5489_out0;
wire v_CARRY_5490_out0;
wire v_CARRY_5491_out0;
wire v_CARRY_5492_out0;
wire v_CARRY_5493_out0;
wire v_CARRY_5494_out0;
wire v_CARRY_5495_out0;
wire v_CARRY_5496_out0;
wire v_CARRY_5497_out0;
wire v_CARRY_5498_out0;
wire v_CARRY_5499_out0;
wire v_CARRY_5500_out0;
wire v_CARRY_5501_out0;
wire v_CARRY_5502_out0;
wire v_CARRY_5503_out0;
wire v_CARRY_5504_out0;
wire v_CARRY_5505_out0;
wire v_CARRY_5506_out0;
wire v_CARRY_5507_out0;
wire v_CARRY_5508_out0;
wire v_CARRY_5509_out0;
wire v_CARRY_5510_out0;
wire v_CARRY_5511_out0;
wire v_CARRY_5512_out0;
wire v_CARRY_5513_out0;
wire v_CARRY_5514_out0;
wire v_CARRY_5515_out0;
wire v_CARRY_5516_out0;
wire v_CARRY_5517_out0;
wire v_CARRY_5518_out0;
wire v_CARRY_5519_out0;
wire v_CARRY_5520_out0;
wire v_CARRY_5521_out0;
wire v_CARRY_5522_out0;
wire v_CARRY_5523_out0;
wire v_CARRY_5524_out0;
wire v_CARRY_5525_out0;
wire v_CARRY_5526_out0;
wire v_CARRY_5527_out0;
wire v_CARRY_5528_out0;
wire v_CARRY_5529_out0;
wire v_CARRY_5530_out0;
wire v_CARRY_5531_out0;
wire v_CARRY_5532_out0;
wire v_CARRY_5533_out0;
wire v_CARRY_5534_out0;
wire v_CARRY_5535_out0;
wire v_CARRY_5536_out0;
wire v_CARRY_5537_out0;
wire v_CARRY_5538_out0;
wire v_CARRY_5539_out0;
wire v_CARRY_5540_out0;
wire v_CARRY_5541_out0;
wire v_CARRY_5542_out0;
wire v_CARRY_5543_out0;
wire v_CARRY_5544_out0;
wire v_CARRY_5545_out0;
wire v_CARRY_5546_out0;
wire v_CARRY_5547_out0;
wire v_CARRY_5548_out0;
wire v_CARRY_5549_out0;
wire v_CARRY_5550_out0;
wire v_CARRY_5551_out0;
wire v_CARRY_5552_out0;
wire v_CARRY_5553_out0;
wire v_CARRY_5554_out0;
wire v_CARRY_5555_out0;
wire v_CARRY_5556_out0;
wire v_CARRY_5557_out0;
wire v_CARRY_5558_out0;
wire v_CARRY_5559_out0;
wire v_CARRY_5560_out0;
wire v_CARRY_5561_out0;
wire v_CARRY_5562_out0;
wire v_CARRY_5563_out0;
wire v_CARRY_5564_out0;
wire v_CARRY_5565_out0;
wire v_CARRY_5566_out0;
wire v_CARRY_5567_out0;
wire v_CARRY_5568_out0;
wire v_CARRY_5569_out0;
wire v_CARRY_5570_out0;
wire v_CARRY_5571_out0;
wire v_CARRY_5572_out0;
wire v_CARRY_5573_out0;
wire v_CARRY_5574_out0;
wire v_CARRY_5575_out0;
wire v_CARRY_5576_out0;
wire v_CARRY_5577_out0;
wire v_CARRY_5578_out0;
wire v_CARRY_5579_out0;
wire v_CARRY_5580_out0;
wire v_CARRY_5581_out0;
wire v_CARRY_5582_out0;
wire v_CARRY_5583_out0;
wire v_CARRY_5584_out0;
wire v_CARRY_5585_out0;
wire v_CARRY_5586_out0;
wire v_CARRY_5587_out0;
wire v_CARRY_5588_out0;
wire v_CARRY_5589_out0;
wire v_CARRY_5590_out0;
wire v_CARRY_5591_out0;
wire v_CARRY_5592_out0;
wire v_CARRY_5593_out0;
wire v_CARRY_5594_out0;
wire v_CARRY_5595_out0;
wire v_CARRY_5596_out0;
wire v_CARRY_5597_out0;
wire v_CARRY_5598_out0;
wire v_CARRY_5599_out0;
wire v_CARRY_5600_out0;
wire v_CARRY_5601_out0;
wire v_CARRY_5602_out0;
wire v_CARRY_5603_out0;
wire v_CARRY_5604_out0;
wire v_CARRY_5605_out0;
wire v_CARRY_5606_out0;
wire v_CARRY_5607_out0;
wire v_CARRY_5608_out0;
wire v_CARRY_5609_out0;
wire v_CARRY_5610_out0;
wire v_CARRY_5611_out0;
wire v_CARRY_5612_out0;
wire v_CARRY_5613_out0;
wire v_CARRY_5614_out0;
wire v_CARRY_5615_out0;
wire v_CARRY_5616_out0;
wire v_CARRY_5617_out0;
wire v_CARRY_5618_out0;
wire v_CARRY_5619_out0;
wire v_CARRY_5620_out0;
wire v_CARRY_5621_out0;
wire v_CARRY_5622_out0;
wire v_CARRY_5623_out0;
wire v_CARRY_5624_out0;
wire v_CARRY_5625_out0;
wire v_CARRY_5626_out0;
wire v_CARRY_5627_out0;
wire v_CARRY_5628_out0;
wire v_CARRY_5629_out0;
wire v_CARRY_5630_out0;
wire v_CARRY_5631_out0;
wire v_CARRY_5632_out0;
wire v_CARRY_5633_out0;
wire v_CARRY_5634_out0;
wire v_CARRY_5635_out0;
wire v_CARRY_5636_out0;
wire v_CARRY_5637_out0;
wire v_CARRY_5638_out0;
wire v_CARRY_5639_out0;
wire v_CARRY_5640_out0;
wire v_CARRY_5641_out0;
wire v_CARRY_5642_out0;
wire v_CARRY_5643_out0;
wire v_CARRY_5644_out0;
wire v_CARRY_5645_out0;
wire v_CARRY_5646_out0;
wire v_CARRY_5647_out0;
wire v_CARRY_5648_out0;
wire v_CARRY_5649_out0;
wire v_CARRY_5650_out0;
wire v_CARRY_5651_out0;
wire v_CARRY_5652_out0;
wire v_CARRY_5653_out0;
wire v_CARRY_5654_out0;
wire v_CARRY_5655_out0;
wire v_CARRY_5656_out0;
wire v_CARRY_5657_out0;
wire v_CARRY_5658_out0;
wire v_CARRY_5659_out0;
wire v_CARRY_5660_out0;
wire v_CARRY_5661_out0;
wire v_CARRY_5662_out0;
wire v_CARRY_5663_out0;
wire v_CARRY_5664_out0;
wire v_CARRY_5665_out0;
wire v_CARRY_5666_out0;
wire v_CARRY_5667_out0;
wire v_CARRY_5668_out0;
wire v_CARRY_5669_out0;
wire v_CARRY_5670_out0;
wire v_CARRY_5671_out0;
wire v_CARRY_5672_out0;
wire v_CARRY_5673_out0;
wire v_CARRY_5674_out0;
wire v_CARRY_5675_out0;
wire v_CARRY_5676_out0;
wire v_CARRY_5677_out0;
wire v_CARRY_5678_out0;
wire v_CARRY_5679_out0;
wire v_CARRY_5680_out0;
wire v_CARRY_5681_out0;
wire v_CARRY_5682_out0;
wire v_CARRY_5683_out0;
wire v_CARRY_5684_out0;
wire v_CARRY_5685_out0;
wire v_CARRY_5686_out0;
wire v_CARRY_5687_out0;
wire v_CARRY_5688_out0;
wire v_CARRY_5689_out0;
wire v_CARRY_5690_out0;
wire v_CARRY_5691_out0;
wire v_CARRY_5692_out0;
wire v_CARRY_5693_out0;
wire v_CARRY_5694_out0;
wire v_CARRY_5695_out0;
wire v_CARRY_5696_out0;
wire v_CARRY_5697_out0;
wire v_CARRY_5698_out0;
wire v_CARRY_5699_out0;
wire v_CARRY_5700_out0;
wire v_CARRY_5701_out0;
wire v_CARRY_5702_out0;
wire v_CARRY_5703_out0;
wire v_CARRY_5704_out0;
wire v_CARRY_5705_out0;
wire v_CARRY_5706_out0;
wire v_CARRY_5707_out0;
wire v_CARRY_5708_out0;
wire v_CARRY_5709_out0;
wire v_CARRY_5710_out0;
wire v_CARRY_5711_out0;
wire v_CARRY_5712_out0;
wire v_CARRY_5713_out0;
wire v_CARRY_5714_out0;
wire v_CARRY_5715_out0;
wire v_CARRY_5716_out0;
wire v_CARRY_5717_out0;
wire v_CARRY_5718_out0;
wire v_CARRY_5719_out0;
wire v_CARRY_5720_out0;
wire v_CARRY_5721_out0;
wire v_CARRY_5722_out0;
wire v_CARRY_5723_out0;
wire v_CARRY_5724_out0;
wire v_CARRY_5725_out0;
wire v_CARRY_5726_out0;
wire v_CARRY_5727_out0;
wire v_CARRY_5728_out0;
wire v_CARRY_5729_out0;
wire v_CARRY_5730_out0;
wire v_CARRY_5731_out0;
wire v_CARRY_5732_out0;
wire v_CARRY_5733_out0;
wire v_CARRY_5734_out0;
wire v_CARRY_5735_out0;
wire v_CARRY_5736_out0;
wire v_CARRY_5737_out0;
wire v_CARRY_5738_out0;
wire v_CARRY_5739_out0;
wire v_CARRY_5740_out0;
wire v_CARRY_5741_out0;
wire v_CARRY_5742_out0;
wire v_CARRY_5743_out0;
wire v_CARRY_5744_out0;
wire v_CARRY_5745_out0;
wire v_CARRY_5746_out0;
wire v_CARRY_5747_out0;
wire v_CARRY_5748_out0;
wire v_CARRY_5749_out0;
wire v_CARRY_5750_out0;
wire v_CARRY_5751_out0;
wire v_CARRY_5752_out0;
wire v_CARRY_5753_out0;
wire v_CARRY_5754_out0;
wire v_CARRY_5755_out0;
wire v_CARRY_5756_out0;
wire v_CARRY_5757_out0;
wire v_CARRY_5758_out0;
wire v_CARRY_5759_out0;
wire v_CARRY_5760_out0;
wire v_CARRY_5761_out0;
wire v_CARRY_5762_out0;
wire v_CARRY_5763_out0;
wire v_CARRY_5764_out0;
wire v_CARRY_5765_out0;
wire v_CARRY_5766_out0;
wire v_CARRY_5767_out0;
wire v_CARRY_5768_out0;
wire v_CARRY_5769_out0;
wire v_CARRY_5770_out0;
wire v_CARRY_5771_out0;
wire v_CARRY_5772_out0;
wire v_CARRY_5773_out0;
wire v_CARRY_5774_out0;
wire v_CARRY_5775_out0;
wire v_CARRY_5776_out0;
wire v_CARRY_5777_out0;
wire v_CARRY_5778_out0;
wire v_CARRY_5779_out0;
wire v_CARRY_5780_out0;
wire v_CARRY_5781_out0;
wire v_CARRY_5782_out0;
wire v_CARRY_5783_out0;
wire v_CARRY_5784_out0;
wire v_CARRY_5785_out0;
wire v_CARRY_5786_out0;
wire v_CARRY_5787_out0;
wire v_CARRY_5788_out0;
wire v_CARRY_5789_out0;
wire v_CIN_10000_out0;
wire v_CIN_10001_out0;
wire v_CIN_10002_out0;
wire v_CIN_10003_out0;
wire v_CIN_10004_out0;
wire v_CIN_10005_out0;
wire v_CIN_10006_out0;
wire v_CIN_10007_out0;
wire v_CIN_10008_out0;
wire v_CIN_10009_out0;
wire v_CIN_10010_out0;
wire v_CIN_10011_out0;
wire v_CIN_10012_out0;
wire v_CIN_10013_out0;
wire v_CIN_10014_out0;
wire v_CIN_10015_out0;
wire v_CIN_10016_out0;
wire v_CIN_10017_out0;
wire v_CIN_10018_out0;
wire v_CIN_10019_out0;
wire v_CIN_10020_out0;
wire v_CIN_10021_out0;
wire v_CIN_10022_out0;
wire v_CIN_10023_out0;
wire v_CIN_10024_out0;
wire v_CIN_10025_out0;
wire v_CIN_10026_out0;
wire v_CIN_10027_out0;
wire v_CIN_10028_out0;
wire v_CIN_10029_out0;
wire v_CIN_10030_out0;
wire v_CIN_10031_out0;
wire v_CIN_10032_out0;
wire v_CIN_10033_out0;
wire v_CIN_10034_out0;
wire v_CIN_10035_out0;
wire v_CIN_10036_out0;
wire v_CIN_10037_out0;
wire v_CIN_10038_out0;
wire v_CIN_10039_out0;
wire v_CIN_10040_out0;
wire v_CIN_10041_out0;
wire v_CIN_10042_out0;
wire v_CIN_10043_out0;
wire v_CIN_10044_out0;
wire v_CIN_10045_out0;
wire v_CIN_10046_out0;
wire v_CIN_10047_out0;
wire v_CIN_10048_out0;
wire v_CIN_10049_out0;
wire v_CIN_10050_out0;
wire v_CIN_10051_out0;
wire v_CIN_10052_out0;
wire v_CIN_10053_out0;
wire v_CIN_10054_out0;
wire v_CIN_10055_out0;
wire v_CIN_10056_out0;
wire v_CIN_10057_out0;
wire v_CIN_10058_out0;
wire v_CIN_10059_out0;
wire v_CIN_10060_out0;
wire v_CIN_10061_out0;
wire v_CIN_10062_out0;
wire v_CIN_10063_out0;
wire v_CIN_10064_out0;
wire v_CIN_10065_out0;
wire v_CIN_10066_out0;
wire v_CIN_10067_out0;
wire v_CIN_10068_out0;
wire v_CIN_10069_out0;
wire v_CIN_10070_out0;
wire v_CIN_10071_out0;
wire v_CIN_10072_out0;
wire v_CIN_10073_out0;
wire v_CIN_10074_out0;
wire v_CIN_10075_out0;
wire v_CIN_10076_out0;
wire v_CIN_10077_out0;
wire v_CIN_10078_out0;
wire v_CIN_10079_out0;
wire v_CIN_10080_out0;
wire v_CIN_10081_out0;
wire v_CIN_10082_out0;
wire v_CIN_10083_out0;
wire v_CIN_10084_out0;
wire v_CIN_10085_out0;
wire v_CIN_10086_out0;
wire v_CIN_10087_out0;
wire v_CIN_10088_out0;
wire v_CIN_10089_out0;
wire v_CIN_10090_out0;
wire v_CIN_10091_out0;
wire v_CIN_10092_out0;
wire v_CIN_10093_out0;
wire v_CIN_10094_out0;
wire v_CIN_10095_out0;
wire v_CIN_10096_out0;
wire v_CIN_10097_out0;
wire v_CIN_10098_out0;
wire v_CIN_10099_out0;
wire v_CIN_10100_out0;
wire v_CIN_10101_out0;
wire v_CIN_10102_out0;
wire v_CIN_10103_out0;
wire v_CIN_10104_out0;
wire v_CIN_10105_out0;
wire v_CIN_10106_out0;
wire v_CIN_10107_out0;
wire v_CIN_10108_out0;
wire v_CIN_10109_out0;
wire v_CIN_10110_out0;
wire v_CIN_10111_out0;
wire v_CIN_10112_out0;
wire v_CIN_10113_out0;
wire v_CIN_10114_out0;
wire v_CIN_10115_out0;
wire v_CIN_10116_out0;
wire v_CIN_10117_out0;
wire v_CIN_10118_out0;
wire v_CIN_10119_out0;
wire v_CIN_10120_out0;
wire v_CIN_10121_out0;
wire v_CIN_10122_out0;
wire v_CIN_10123_out0;
wire v_CIN_10124_out0;
wire v_CIN_10125_out0;
wire v_CIN_10126_out0;
wire v_CIN_10127_out0;
wire v_CIN_10128_out0;
wire v_CIN_10129_out0;
wire v_CIN_10130_out0;
wire v_CIN_10131_out0;
wire v_CIN_10132_out0;
wire v_CIN_10133_out0;
wire v_CIN_10134_out0;
wire v_CIN_10135_out0;
wire v_CIN_10136_out0;
wire v_CIN_10137_out0;
wire v_CIN_10138_out0;
wire v_CIN_10139_out0;
wire v_CIN_10140_out0;
wire v_CIN_10141_out0;
wire v_CIN_10142_out0;
wire v_CIN_10143_out0;
wire v_CIN_10144_out0;
wire v_CIN_10145_out0;
wire v_CIN_10146_out0;
wire v_CIN_10147_out0;
wire v_CIN_10148_out0;
wire v_CIN_10149_out0;
wire v_CIN_10150_out0;
wire v_CIN_10151_out0;
wire v_CIN_10152_out0;
wire v_CIN_10153_out0;
wire v_CIN_10154_out0;
wire v_CIN_10155_out0;
wire v_CIN_10156_out0;
wire v_CIN_10157_out0;
wire v_CIN_10158_out0;
wire v_CIN_10159_out0;
wire v_CIN_10160_out0;
wire v_CIN_10161_out0;
wire v_CIN_10162_out0;
wire v_CIN_10163_out0;
wire v_CIN_10164_out0;
wire v_CIN_10165_out0;
wire v_CIN_10166_out0;
wire v_CIN_10167_out0;
wire v_CIN_10168_out0;
wire v_CIN_10169_out0;
wire v_CIN_10170_out0;
wire v_CIN_10171_out0;
wire v_CIN_10172_out0;
wire v_CIN_10173_out0;
wire v_CIN_10174_out0;
wire v_CIN_10175_out0;
wire v_CIN_10176_out0;
wire v_CIN_10177_out0;
wire v_CIN_10178_out0;
wire v_CIN_10179_out0;
wire v_CIN_10180_out0;
wire v_CIN_10181_out0;
wire v_CIN_10182_out0;
wire v_CIN_10183_out0;
wire v_CIN_10184_out0;
wire v_CIN_10185_out0;
wire v_CIN_10186_out0;
wire v_CIN_10187_out0;
wire v_CIN_10188_out0;
wire v_CIN_10189_out0;
wire v_CIN_10190_out0;
wire v_CIN_10191_out0;
wire v_CIN_10192_out0;
wire v_CIN_10193_out0;
wire v_CIN_10194_out0;
wire v_CIN_10195_out0;
wire v_CIN_10196_out0;
wire v_CIN_10197_out0;
wire v_CIN_10198_out0;
wire v_CIN_10199_out0;
wire v_CIN_10200_out0;
wire v_CIN_10201_out0;
wire v_CIN_10202_out0;
wire v_CIN_10203_out0;
wire v_CIN_10204_out0;
wire v_CIN_10205_out0;
wire v_CIN_10206_out0;
wire v_CIN_10207_out0;
wire v_CIN_10208_out0;
wire v_CIN_10209_out0;
wire v_CIN_10210_out0;
wire v_CIN_10211_out0;
wire v_CIN_10212_out0;
wire v_CIN_10213_out0;
wire v_CIN_10214_out0;
wire v_CIN_10215_out0;
wire v_CIN_10216_out0;
wire v_CIN_10217_out0;
wire v_CIN_10218_out0;
wire v_CIN_10219_out0;
wire v_CIN_10220_out0;
wire v_CIN_10221_out0;
wire v_CIN_10222_out0;
wire v_CIN_10223_out0;
wire v_CIN_10224_out0;
wire v_CIN_10225_out0;
wire v_CIN_10226_out0;
wire v_CIN_10227_out0;
wire v_CIN_10228_out0;
wire v_CIN_10229_out0;
wire v_CIN_10230_out0;
wire v_CIN_10231_out0;
wire v_CIN_10232_out0;
wire v_CIN_10233_out0;
wire v_CIN_10234_out0;
wire v_CIN_10235_out0;
wire v_CIN_10236_out0;
wire v_CIN_10237_out0;
wire v_CIN_10238_out0;
wire v_CIN_10239_out0;
wire v_CIN_10240_out0;
wire v_CIN_10241_out0;
wire v_CIN_10242_out0;
wire v_CIN_10243_out0;
wire v_CIN_10244_out0;
wire v_CIN_10245_out0;
wire v_CIN_10246_out0;
wire v_CIN_10247_out0;
wire v_CIN_10248_out0;
wire v_CIN_10249_out0;
wire v_CIN_10250_out0;
wire v_CIN_10251_out0;
wire v_CIN_10252_out0;
wire v_CIN_10253_out0;
wire v_CIN_10254_out0;
wire v_CIN_10255_out0;
wire v_CIN_9808_out0;
wire v_CIN_9809_out0;
wire v_CIN_9810_out0;
wire v_CIN_9811_out0;
wire v_CIN_9812_out0;
wire v_CIN_9813_out0;
wire v_CIN_9814_out0;
wire v_CIN_9815_out0;
wire v_CIN_9816_out0;
wire v_CIN_9817_out0;
wire v_CIN_9818_out0;
wire v_CIN_9819_out0;
wire v_CIN_9820_out0;
wire v_CIN_9821_out0;
wire v_CIN_9822_out0;
wire v_CIN_9823_out0;
wire v_CIN_9824_out0;
wire v_CIN_9825_out0;
wire v_CIN_9826_out0;
wire v_CIN_9827_out0;
wire v_CIN_9828_out0;
wire v_CIN_9829_out0;
wire v_CIN_9830_out0;
wire v_CIN_9831_out0;
wire v_CIN_9832_out0;
wire v_CIN_9833_out0;
wire v_CIN_9834_out0;
wire v_CIN_9835_out0;
wire v_CIN_9836_out0;
wire v_CIN_9837_out0;
wire v_CIN_9838_out0;
wire v_CIN_9839_out0;
wire v_CIN_9840_out0;
wire v_CIN_9841_out0;
wire v_CIN_9842_out0;
wire v_CIN_9843_out0;
wire v_CIN_9844_out0;
wire v_CIN_9845_out0;
wire v_CIN_9846_out0;
wire v_CIN_9847_out0;
wire v_CIN_9848_out0;
wire v_CIN_9849_out0;
wire v_CIN_9850_out0;
wire v_CIN_9851_out0;
wire v_CIN_9852_out0;
wire v_CIN_9853_out0;
wire v_CIN_9854_out0;
wire v_CIN_9855_out0;
wire v_CIN_9856_out0;
wire v_CIN_9857_out0;
wire v_CIN_9858_out0;
wire v_CIN_9859_out0;
wire v_CIN_9860_out0;
wire v_CIN_9861_out0;
wire v_CIN_9862_out0;
wire v_CIN_9863_out0;
wire v_CIN_9864_out0;
wire v_CIN_9865_out0;
wire v_CIN_9866_out0;
wire v_CIN_9867_out0;
wire v_CIN_9868_out0;
wire v_CIN_9869_out0;
wire v_CIN_9870_out0;
wire v_CIN_9871_out0;
wire v_CIN_9872_out0;
wire v_CIN_9873_out0;
wire v_CIN_9874_out0;
wire v_CIN_9875_out0;
wire v_CIN_9876_out0;
wire v_CIN_9877_out0;
wire v_CIN_9878_out0;
wire v_CIN_9879_out0;
wire v_CIN_9880_out0;
wire v_CIN_9881_out0;
wire v_CIN_9882_out0;
wire v_CIN_9883_out0;
wire v_CIN_9884_out0;
wire v_CIN_9885_out0;
wire v_CIN_9886_out0;
wire v_CIN_9887_out0;
wire v_CIN_9888_out0;
wire v_CIN_9889_out0;
wire v_CIN_9890_out0;
wire v_CIN_9891_out0;
wire v_CIN_9892_out0;
wire v_CIN_9893_out0;
wire v_CIN_9894_out0;
wire v_CIN_9895_out0;
wire v_CIN_9896_out0;
wire v_CIN_9897_out0;
wire v_CIN_9898_out0;
wire v_CIN_9899_out0;
wire v_CIN_9900_out0;
wire v_CIN_9901_out0;
wire v_CIN_9902_out0;
wire v_CIN_9903_out0;
wire v_CIN_9904_out0;
wire v_CIN_9905_out0;
wire v_CIN_9906_out0;
wire v_CIN_9907_out0;
wire v_CIN_9908_out0;
wire v_CIN_9909_out0;
wire v_CIN_9910_out0;
wire v_CIN_9911_out0;
wire v_CIN_9912_out0;
wire v_CIN_9913_out0;
wire v_CIN_9914_out0;
wire v_CIN_9915_out0;
wire v_CIN_9916_out0;
wire v_CIN_9917_out0;
wire v_CIN_9918_out0;
wire v_CIN_9919_out0;
wire v_CIN_9920_out0;
wire v_CIN_9921_out0;
wire v_CIN_9922_out0;
wire v_CIN_9923_out0;
wire v_CIN_9924_out0;
wire v_CIN_9925_out0;
wire v_CIN_9926_out0;
wire v_CIN_9927_out0;
wire v_CIN_9928_out0;
wire v_CIN_9929_out0;
wire v_CIN_9930_out0;
wire v_CIN_9931_out0;
wire v_CIN_9932_out0;
wire v_CIN_9933_out0;
wire v_CIN_9934_out0;
wire v_CIN_9935_out0;
wire v_CIN_9936_out0;
wire v_CIN_9937_out0;
wire v_CIN_9938_out0;
wire v_CIN_9939_out0;
wire v_CIN_9940_out0;
wire v_CIN_9941_out0;
wire v_CIN_9942_out0;
wire v_CIN_9943_out0;
wire v_CIN_9944_out0;
wire v_CIN_9945_out0;
wire v_CIN_9946_out0;
wire v_CIN_9947_out0;
wire v_CIN_9948_out0;
wire v_CIN_9949_out0;
wire v_CIN_9950_out0;
wire v_CIN_9951_out0;
wire v_CIN_9952_out0;
wire v_CIN_9953_out0;
wire v_CIN_9954_out0;
wire v_CIN_9955_out0;
wire v_CIN_9956_out0;
wire v_CIN_9957_out0;
wire v_CIN_9958_out0;
wire v_CIN_9959_out0;
wire v_CIN_9960_out0;
wire v_CIN_9961_out0;
wire v_CIN_9962_out0;
wire v_CIN_9963_out0;
wire v_CIN_9964_out0;
wire v_CIN_9965_out0;
wire v_CIN_9966_out0;
wire v_CIN_9967_out0;
wire v_CIN_9968_out0;
wire v_CIN_9969_out0;
wire v_CIN_9970_out0;
wire v_CIN_9971_out0;
wire v_CIN_9972_out0;
wire v_CIN_9973_out0;
wire v_CIN_9974_out0;
wire v_CIN_9975_out0;
wire v_CIN_9976_out0;
wire v_CIN_9977_out0;
wire v_CIN_9978_out0;
wire v_CIN_9979_out0;
wire v_CIN_9980_out0;
wire v_CIN_9981_out0;
wire v_CIN_9982_out0;
wire v_CIN_9983_out0;
wire v_CIN_9984_out0;
wire v_CIN_9985_out0;
wire v_CIN_9986_out0;
wire v_CIN_9987_out0;
wire v_CIN_9988_out0;
wire v_CIN_9989_out0;
wire v_CIN_9990_out0;
wire v_CIN_9991_out0;
wire v_CIN_9992_out0;
wire v_CIN_9993_out0;
wire v_CIN_9994_out0;
wire v_CIN_9995_out0;
wire v_CIN_9996_out0;
wire v_CIN_9997_out0;
wire v_CIN_9998_out0;
wire v_CIN_9999_out0;
wire v_CMP_13609_out0;
wire v_CMP_13610_out0;
wire v_CMP_3805_out0;
wire v_CMP_3806_out0;
wire v_CMP_8646_out0;
wire v_CMP_8647_out0;
wire v_COUT_1000_out0;
wire v_COUT_1001_out0;
wire v_COUT_1002_out0;
wire v_COUT_1003_out0;
wire v_COUT_1004_out0;
wire v_COUT_1005_out0;
wire v_COUT_1006_out0;
wire v_COUT_1007_out0;
wire v_COUT_1008_out0;
wire v_COUT_1009_out0;
wire v_COUT_1010_out0;
wire v_COUT_1011_out0;
wire v_COUT_1012_out0;
wire v_COUT_1013_out0;
wire v_COUT_1014_out0;
wire v_COUT_1015_out0;
wire v_COUT_1016_out0;
wire v_COUT_1017_out0;
wire v_COUT_1018_out0;
wire v_COUT_1019_out0;
wire v_COUT_1020_out0;
wire v_COUT_1021_out0;
wire v_COUT_1022_out0;
wire v_COUT_1023_out0;
wire v_COUT_1024_out0;
wire v_COUT_1025_out0;
wire v_COUT_1026_out0;
wire v_COUT_1027_out0;
wire v_COUT_1028_out0;
wire v_COUT_1029_out0;
wire v_COUT_1030_out0;
wire v_COUT_1031_out0;
wire v_COUT_1032_out0;
wire v_COUT_1033_out0;
wire v_COUT_1034_out0;
wire v_COUT_1035_out0;
wire v_COUT_1036_out0;
wire v_COUT_1037_out0;
wire v_COUT_1038_out0;
wire v_COUT_1039_out0;
wire v_COUT_1040_out0;
wire v_COUT_1041_out0;
wire v_COUT_1042_out0;
wire v_COUT_1043_out0;
wire v_COUT_1044_out0;
wire v_COUT_1045_out0;
wire v_COUT_1046_out0;
wire v_COUT_1047_out0;
wire v_COUT_1048_out0;
wire v_COUT_1049_out0;
wire v_COUT_1050_out0;
wire v_COUT_1051_out0;
wire v_COUT_1052_out0;
wire v_COUT_1053_out0;
wire v_COUT_10547_out0;
wire v_COUT_10548_out0;
wire v_COUT_1054_out0;
wire v_COUT_1055_out0;
wire v_COUT_1056_out0;
wire v_COUT_1057_out0;
wire v_COUT_1058_out0;
wire v_COUT_1059_out0;
wire v_COUT_1060_out0;
wire v_COUT_1061_out0;
wire v_COUT_1062_out0;
wire v_COUT_1063_out0;
wire v_COUT_1064_out0;
wire v_COUT_1065_out0;
wire v_COUT_1066_out0;
wire v_COUT_1067_out0;
wire v_COUT_1068_out0;
wire v_COUT_1069_out0;
wire v_COUT_1070_out0;
wire v_COUT_1071_out0;
wire v_COUT_1072_out0;
wire v_COUT_1073_out0;
wire v_COUT_1074_out0;
wire v_COUT_1075_out0;
wire v_COUT_1076_out0;
wire v_COUT_1077_out0;
wire v_COUT_1078_out0;
wire v_COUT_1079_out0;
wire v_COUT_1080_out0;
wire v_COUT_1081_out0;
wire v_COUT_1082_out0;
wire v_COUT_1083_out0;
wire v_COUT_1084_out0;
wire v_COUT_1085_out0;
wire v_COUT_1086_out0;
wire v_COUT_1087_out0;
wire v_COUT_1088_out0;
wire v_COUT_1089_out0;
wire v_COUT_1090_out0;
wire v_COUT_1091_out0;
wire v_COUT_1092_out0;
wire v_COUT_1093_out0;
wire v_COUT_1094_out0;
wire v_COUT_1095_out0;
wire v_COUT_1096_out0;
wire v_COUT_1097_out0;
wire v_COUT_1098_out0;
wire v_COUT_1099_out0;
wire v_COUT_1100_out0;
wire v_COUT_1101_out0;
wire v_COUT_1102_out0;
wire v_COUT_1103_out0;
wire v_COUT_1104_out0;
wire v_COUT_1105_out0;
wire v_COUT_1106_out0;
wire v_COUT_1107_out0;
wire v_COUT_1108_out0;
wire v_COUT_1109_out0;
wire v_COUT_1110_out0;
wire v_COUT_1111_out0;
wire v_COUT_1112_out0;
wire v_COUT_1113_out0;
wire v_COUT_1114_out0;
wire v_COUT_1115_out0;
wire v_COUT_1116_out0;
wire v_COUT_1117_out0;
wire v_COUT_1118_out0;
wire v_COUT_1119_out0;
wire v_COUT_1120_out0;
wire v_COUT_1121_out0;
wire v_COUT_1122_out0;
wire v_COUT_1123_out0;
wire v_COUT_1124_out0;
wire v_COUT_1125_out0;
wire v_COUT_1126_out0;
wire v_COUT_1127_out0;
wire v_COUT_1128_out0;
wire v_COUT_1129_out0;
wire v_COUT_1130_out0;
wire v_COUT_1131_out0;
wire v_COUT_1132_out0;
wire v_COUT_1133_out0;
wire v_COUT_1134_out0;
wire v_COUT_2725_out0;
wire v_COUT_3895_out0;
wire v_COUT_3896_out0;
wire v_COUT_687_out0;
wire v_COUT_688_out0;
wire v_COUT_689_out0;
wire v_COUT_690_out0;
wire v_COUT_691_out0;
wire v_COUT_692_out0;
wire v_COUT_693_out0;
wire v_COUT_694_out0;
wire v_COUT_695_out0;
wire v_COUT_696_out0;
wire v_COUT_697_out0;
wire v_COUT_698_out0;
wire v_COUT_699_out0;
wire v_COUT_700_out0;
wire v_COUT_701_out0;
wire v_COUT_702_out0;
wire v_COUT_703_out0;
wire v_COUT_704_out0;
wire v_COUT_705_out0;
wire v_COUT_706_out0;
wire v_COUT_707_out0;
wire v_COUT_708_out0;
wire v_COUT_709_out0;
wire v_COUT_70_out0;
wire v_COUT_710_out0;
wire v_COUT_711_out0;
wire v_COUT_712_out0;
wire v_COUT_713_out0;
wire v_COUT_714_out0;
wire v_COUT_715_out0;
wire v_COUT_716_out0;
wire v_COUT_717_out0;
wire v_COUT_718_out0;
wire v_COUT_719_out0;
wire v_COUT_71_out0;
wire v_COUT_720_out0;
wire v_COUT_721_out0;
wire v_COUT_722_out0;
wire v_COUT_723_out0;
wire v_COUT_724_out0;
wire v_COUT_725_out0;
wire v_COUT_726_out0;
wire v_COUT_727_out0;
wire v_COUT_728_out0;
wire v_COUT_729_out0;
wire v_COUT_730_out0;
wire v_COUT_731_out0;
wire v_COUT_732_out0;
wire v_COUT_733_out0;
wire v_COUT_734_out0;
wire v_COUT_735_out0;
wire v_COUT_736_out0;
wire v_COUT_737_out0;
wire v_COUT_738_out0;
wire v_COUT_739_out0;
wire v_COUT_740_out0;
wire v_COUT_741_out0;
wire v_COUT_742_out0;
wire v_COUT_743_out0;
wire v_COUT_744_out0;
wire v_COUT_745_out0;
wire v_COUT_746_out0;
wire v_COUT_747_out0;
wire v_COUT_748_out0;
wire v_COUT_749_out0;
wire v_COUT_750_out0;
wire v_COUT_751_out0;
wire v_COUT_752_out0;
wire v_COUT_753_out0;
wire v_COUT_754_out0;
wire v_COUT_755_out0;
wire v_COUT_756_out0;
wire v_COUT_757_out0;
wire v_COUT_758_out0;
wire v_COUT_759_out0;
wire v_COUT_760_out0;
wire v_COUT_761_out0;
wire v_COUT_762_out0;
wire v_COUT_763_out0;
wire v_COUT_764_out0;
wire v_COUT_765_out0;
wire v_COUT_766_out0;
wire v_COUT_767_out0;
wire v_COUT_768_out0;
wire v_COUT_769_out0;
wire v_COUT_770_out0;
wire v_COUT_771_out0;
wire v_COUT_772_out0;
wire v_COUT_773_out0;
wire v_COUT_774_out0;
wire v_COUT_775_out0;
wire v_COUT_776_out0;
wire v_COUT_777_out0;
wire v_COUT_778_out0;
wire v_COUT_779_out0;
wire v_COUT_780_out0;
wire v_COUT_781_out0;
wire v_COUT_782_out0;
wire v_COUT_783_out0;
wire v_COUT_784_out0;
wire v_COUT_785_out0;
wire v_COUT_786_out0;
wire v_COUT_787_out0;
wire v_COUT_788_out0;
wire v_COUT_789_out0;
wire v_COUT_790_out0;
wire v_COUT_791_out0;
wire v_COUT_792_out0;
wire v_COUT_793_out0;
wire v_COUT_794_out0;
wire v_COUT_795_out0;
wire v_COUT_796_out0;
wire v_COUT_797_out0;
wire v_COUT_798_out0;
wire v_COUT_799_out0;
wire v_COUT_800_out0;
wire v_COUT_801_out0;
wire v_COUT_802_out0;
wire v_COUT_803_out0;
wire v_COUT_804_out0;
wire v_COUT_805_out0;
wire v_COUT_806_out0;
wire v_COUT_807_out0;
wire v_COUT_808_out0;
wire v_COUT_809_out0;
wire v_COUT_810_out0;
wire v_COUT_811_out0;
wire v_COUT_812_out0;
wire v_COUT_813_out0;
wire v_COUT_814_out0;
wire v_COUT_815_out0;
wire v_COUT_816_out0;
wire v_COUT_817_out0;
wire v_COUT_818_out0;
wire v_COUT_819_out0;
wire v_COUT_820_out0;
wire v_COUT_821_out0;
wire v_COUT_822_out0;
wire v_COUT_823_out0;
wire v_COUT_824_out0;
wire v_COUT_825_out0;
wire v_COUT_826_out0;
wire v_COUT_827_out0;
wire v_COUT_828_out0;
wire v_COUT_829_out0;
wire v_COUT_830_out0;
wire v_COUT_831_out0;
wire v_COUT_832_out0;
wire v_COUT_833_out0;
wire v_COUT_834_out0;
wire v_COUT_835_out0;
wire v_COUT_836_out0;
wire v_COUT_837_out0;
wire v_COUT_838_out0;
wire v_COUT_839_out0;
wire v_COUT_840_out0;
wire v_COUT_841_out0;
wire v_COUT_842_out0;
wire v_COUT_843_out0;
wire v_COUT_844_out0;
wire v_COUT_845_out0;
wire v_COUT_846_out0;
wire v_COUT_847_out0;
wire v_COUT_848_out0;
wire v_COUT_849_out0;
wire v_COUT_850_out0;
wire v_COUT_851_out0;
wire v_COUT_852_out0;
wire v_COUT_853_out0;
wire v_COUT_854_out0;
wire v_COUT_855_out0;
wire v_COUT_856_out0;
wire v_COUT_857_out0;
wire v_COUT_858_out0;
wire v_COUT_859_out0;
wire v_COUT_860_out0;
wire v_COUT_861_out0;
wire v_COUT_862_out0;
wire v_COUT_863_out0;
wire v_COUT_864_out0;
wire v_COUT_865_out0;
wire v_COUT_866_out0;
wire v_COUT_867_out0;
wire v_COUT_868_out0;
wire v_COUT_869_out0;
wire v_COUT_870_out0;
wire v_COUT_871_out0;
wire v_COUT_872_out0;
wire v_COUT_873_out0;
wire v_COUT_874_out0;
wire v_COUT_875_out0;
wire v_COUT_876_out0;
wire v_COUT_877_out0;
wire v_COUT_878_out0;
wire v_COUT_879_out0;
wire v_COUT_880_out0;
wire v_COUT_881_out0;
wire v_COUT_882_out0;
wire v_COUT_883_out0;
wire v_COUT_884_out0;
wire v_COUT_885_out0;
wire v_COUT_886_out0;
wire v_COUT_887_out0;
wire v_COUT_888_out0;
wire v_COUT_889_out0;
wire v_COUT_890_out0;
wire v_COUT_891_out0;
wire v_COUT_892_out0;
wire v_COUT_893_out0;
wire v_COUT_894_out0;
wire v_COUT_895_out0;
wire v_COUT_896_out0;
wire v_COUT_897_out0;
wire v_COUT_898_out0;
wire v_COUT_899_out0;
wire v_COUT_900_out0;
wire v_COUT_901_out0;
wire v_COUT_902_out0;
wire v_COUT_903_out0;
wire v_COUT_904_out0;
wire v_COUT_905_out0;
wire v_COUT_906_out0;
wire v_COUT_907_out0;
wire v_COUT_908_out0;
wire v_COUT_909_out0;
wire v_COUT_910_out0;
wire v_COUT_911_out0;
wire v_COUT_912_out0;
wire v_COUT_913_out0;
wire v_COUT_914_out0;
wire v_COUT_915_out0;
wire v_COUT_916_out0;
wire v_COUT_917_out0;
wire v_COUT_918_out0;
wire v_COUT_919_out0;
wire v_COUT_920_out0;
wire v_COUT_921_out0;
wire v_COUT_922_out0;
wire v_COUT_923_out0;
wire v_COUT_924_out0;
wire v_COUT_925_out0;
wire v_COUT_926_out0;
wire v_COUT_927_out0;
wire v_COUT_928_out0;
wire v_COUT_929_out0;
wire v_COUT_930_out0;
wire v_COUT_931_out0;
wire v_COUT_932_out0;
wire v_COUT_933_out0;
wire v_COUT_934_out0;
wire v_COUT_935_out0;
wire v_COUT_936_out0;
wire v_COUT_937_out0;
wire v_COUT_938_out0;
wire v_COUT_939_out0;
wire v_COUT_940_out0;
wire v_COUT_941_out0;
wire v_COUT_942_out0;
wire v_COUT_943_out0;
wire v_COUT_944_out0;
wire v_COUT_945_out0;
wire v_COUT_946_out0;
wire v_COUT_947_out0;
wire v_COUT_948_out0;
wire v_COUT_949_out0;
wire v_COUT_950_out0;
wire v_COUT_951_out0;
wire v_COUT_952_out0;
wire v_COUT_953_out0;
wire v_COUT_954_out0;
wire v_COUT_955_out0;
wire v_COUT_956_out0;
wire v_COUT_957_out0;
wire v_COUT_958_out0;
wire v_COUT_959_out0;
wire v_COUT_960_out0;
wire v_COUT_961_out0;
wire v_COUT_962_out0;
wire v_COUT_963_out0;
wire v_COUT_964_out0;
wire v_COUT_965_out0;
wire v_COUT_966_out0;
wire v_COUT_967_out0;
wire v_COUT_968_out0;
wire v_COUT_969_out0;
wire v_COUT_970_out0;
wire v_COUT_971_out0;
wire v_COUT_972_out0;
wire v_COUT_973_out0;
wire v_COUT_974_out0;
wire v_COUT_975_out0;
wire v_COUT_976_out0;
wire v_COUT_977_out0;
wire v_COUT_978_out0;
wire v_COUT_979_out0;
wire v_COUT_980_out0;
wire v_COUT_981_out0;
wire v_COUT_982_out0;
wire v_COUT_983_out0;
wire v_COUT_984_out0;
wire v_COUT_985_out0;
wire v_COUT_986_out0;
wire v_COUT_987_out0;
wire v_COUT_988_out0;
wire v_COUT_989_out0;
wire v_COUT_990_out0;
wire v_COUT_991_out0;
wire v_COUT_992_out0;
wire v_COUT_993_out0;
wire v_COUT_994_out0;
wire v_COUT_995_out0;
wire v_COUT_996_out0;
wire v_COUT_997_out0;
wire v_COUT_998_out0;
wire v_COUT_999_out0;
wire v_C_13767_out0;
wire v_C_13768_out0;
wire v_C_238_out0;
wire v_C_239_out0;
wire v_C_3197_out0;
wire v_C_3198_out0;
wire v_C_3207_out0;
wire v_C_3208_out0;
wire v_C_379_out0;
wire v_C_380_out0;
wire v_C_4848_out0;
wire v_C_4849_out0;
wire v_C_8648_out0;
wire v_C_8649_out0;
wire v_C_8653_out0;
wire v_C_8654_out0;
wire v_D1_8842_out0;
wire v_D1_8842_out1;
wire v_D1_8842_out2;
wire v_D1_8842_out3;
wire v_D1_8843_out0;
wire v_D1_8843_out1;
wire v_D1_8843_out2;
wire v_D1_8843_out3;
wire v_DIV_INSTRUCTION_11296_out0;
wire v_DIV_INSTRUCTION_11297_out0;
wire v_DIV_INSTRUCTION_13635_out0;
wire v_DIV_INSTRUCTION_13636_out0;
wire v_DIV_INSTRUCTION_3296_out0;
wire v_DIV_INSTRUCTION_3297_out0;
wire v_DIV_INSTRUCTION_4614_out0;
wire v_DIV_INSTRUCTION_4615_out0;
wire v_DIV_INST_2324_out0;
wire v_DIV_INST_2325_out0;
wire v_DONE_RECEIVING_3084_out0;
wire v_DONE_RECEIVING_5857_out0;
wire v_D_7679_out0;
wire v_D_7680_out0;
wire v_D_7681_out0;
wire v_D_7682_out0;
wire v_D_7683_out0;
wire v_D_7684_out0;
wire v_D_7685_out0;
wire v_D_7686_out0;
wire v_D_7687_out0;
wire v_D_7688_out0;
wire v_D_7689_out0;
wire v_D_7690_out0;
wire v_D_7691_out0;
wire v_D_7692_out0;
wire v_D_7693_out0;
wire v_D_7694_out0;
wire v_ENABLE_1757_out0;
wire v_ENABLE_2018_out0;
wire v_ENABLE_2019_out0;
wire v_ENABLE_2020_out0;
wire v_ENABLE_2021_out0;
wire v_ENABLE_2651_out0;
wire v_EN_10451_out0;
wire v_EN_10452_out0;
wire v_EN_10453_out0;
wire v_EN_10454_out0;
wire v_EN_10474_out0;
wire v_EN_10475_out0;
wire v_EN_13181_out0;
wire v_EN_13182_out0;
wire v_EN_2330_out0;
wire v_EN_2331_out0;
wire v_EN_2445_out0;
wire v_EN_2446_out0;
wire v_EN_2919_out0;
wire v_EN_2920_out0;
wire v_EN_2921_out0;
wire v_EN_2922_out0;
wire v_EN_2923_out0;
wire v_EN_2924_out0;
wire v_EN_2925_out0;
wire v_EN_2926_out0;
wire v_EN_2927_out0;
wire v_EN_2928_out0;
wire v_EN_2929_out0;
wire v_EN_2930_out0;
wire v_EN_2931_out0;
wire v_EN_2932_out0;
wire v_EN_2933_out0;
wire v_EN_2934_out0;
wire v_EN_4485_out0;
wire v_EN_4593_out0;
wire v_EN_4594_out0;
wire v_EN_7093_out0;
wire v_EN_7094_out0;
wire v_EN_STALL_10344_out0;
wire v_EN_STALL_13747_out0;
wire v_EQ01_10510_out0;
wire v_EQ01_10511_out0;
wire v_EQ10_2320_out0;
wire v_EQ10_2321_out0;
wire v_EQ11_2456_out0;
wire v_EQ11_2457_out0;
wire v_EQ11_4465_out0;
wire v_EQ11_4466_out0;
wire v_EQ1_10329_out0;
wire v_EQ1_1157_out0;
wire v_EQ1_1158_out0;
wire v_EQ1_13433_out0;
wire v_EQ1_13434_out0;
wire v_EQ1_1857_out0;
wire v_EQ1_1858_out0;
wire v_EQ1_2540_out0;
wire v_EQ1_2541_out0;
wire v_EQ1_2597_out0;
wire v_EQ1_2598_out0;
wire v_EQ1_2675_out0;
wire v_EQ1_2676_out0;
wire v_EQ1_315_out0;
wire v_EQ1_316_out0;
wire v_EQ1_3344_out0;
wire v_EQ1_6956_out0;
wire v_EQ1_6957_out0;
wire v_EQ1_7098_out0;
wire v_EQ1_7099_out0;
wire v_EQ2_10347_out0;
wire v_EQ2_10348_out0;
wire v_EQ2_10771_out0;
wire v_EQ2_10772_out0;
wire v_EQ2_10981_out0;
wire v_EQ2_11254_out0;
wire v_EQ2_11255_out0;
wire v_EQ2_1753_out0;
wire v_EQ2_1754_out0;
wire v_EQ2_7091_out0;
wire v_EQ2_7092_out0;
wire v_EQ2_8_out0;
wire v_EQ2_9795_out0;
wire v_EQ2_9_out0;
wire v_EQ3_11044_out0;
wire v_EQ3_11045_out0;
wire v_EQ3_13504_out0;
wire v_EQ3_13505_out0;
wire v_EQ3_2966_out0;
wire v_EQ3_2967_out0;
wire v_EQ3_5861_out0;
wire v_EQ3_7126_out0;
wire v_EQ3_7127_out0;
wire v_EQ3_7145_out0;
wire v_EQ3_7146_out0;
wire v_EQ4_10345_out0;
wire v_EQ4_10346_out0;
wire v_EQ4_1142_out0;
wire v_EQ4_2149_out0;
wire v_EQ4_3227_out0;
wire v_EQ4_3228_out0;
wire v_EQ4_611_out0;
wire v_EQ4_612_out0;
wire v_EQ5_10364_out0;
wire v_EQ5_10365_out0;
wire v_EQ5_4860_out0;
wire v_EQ5_4861_out0;
wire v_EQ6_1686_out0;
wire v_EQ6_1687_out0;
wire v_EQ6_1966_out0;
wire v_EQ6_1967_out0;
wire v_EQ6_19_out0;
wire v_EQ6_3257_out0;
wire v_EQ7_10399_out0;
wire v_EQ7_10400_out0;
wire v_EQ7_13769_out0;
wire v_EQ7_3307_out0;
wire v_EQ7_3308_out0;
wire v_EQ8_10804_out0;
wire v_EQ8_10805_out0;
wire v_EQ8_2453_out0;
wire v_EQ8_2454_out0;
wire v_EQ8_2874_out0;
wire v_EQ8_2951_out0;
wire v_EQ8_2952_out0;
wire v_EQ9_2007_out0;
wire v_EQ9_2390_out0;
wire v_EQ9_2391_out0;
wire v_EQ9_4842_out0;
wire v_EQ9_4843_out0;
wire v_EQ_100_out0;
wire v_EQ_101_out0;
wire v_EQ_2591_out0;
wire v_EQ_2592_out0;
wire v_EQ_3821_out0;
wire v_EQ_3822_out0;
wire v_EQ_4835_out0;
wire v_EQ_4836_out0;
wire v_EXEC10_2329_out0;
wire v_EXEC10_8812_out0;
wire v_EXEC11_2830_out0;
wire v_EXEC11_4528_out0;
wire v_EXEC1LS_10506_out0;
wire v_EXEC1LS_10507_out0;
wire v_EXEC1LS_10703_out0;
wire v_EXEC1LS_10704_out0;
wire v_EXEC1LS_10843_out0;
wire v_EXEC1LS_10844_out0;
wire v_EXEC1LS_430_out0;
wire v_EXEC1LS_431_out0;
wire v_EXEC1LS_4697_out0;
wire v_EXEC1LS_4698_out0;
wire v_EXEC1LS_6795_out0;
wire v_EXEC1LS_6796_out0;
wire v_EXEC1_10763_out0;
wire v_EXEC1_10764_out0;
wire v_EXEC1_1863_out0;
wire v_EXEC1_1864_out0;
wire v_EXEC1_20_out0;
wire v_EXEC1_21_out0;
wire v_EXEC1_2634_out0;
wire v_EXEC1_2635_out0;
wire v_EXEC1_3038_out0;
wire v_EXEC1_3039_out0;
wire v_EXEC1_7029_out0;
wire v_EXEC1_7030_out0;
wire v_EXEC1_7128_out0;
wire v_EXEC1_7129_out0;
wire v_EXEC20_629_out0;
wire v_EXEC2LS_10549_out0;
wire v_EXEC2LS_10979_out0;
wire v_EXEC2LS_10980_out0;
wire v_EXEC2LS_13558_out0;
wire v_EXEC2LS_13559_out0;
wire v_EXEC2LS_2844_out0;
wire v_EXEC2LS_2845_out0;
wire v_EXEC2LS_3081_out0;
wire v_EXEC2LS_3082_out0;
wire v_EXEC2LS_3188_out0;
wire v_EXEC2LS_3189_out0;
wire v_EXEC2LS_3231_out0;
wire v_EXEC2LS_3232_out0;
wire v_EXEC2_2010_out0;
wire v_EXEC2_2011_out0;
wire v_EXEC2_2110_out0;
wire v_EXEC2_2111_out0;
wire v_EXEC2_2647_out0;
wire v_EXEC2_2648_out0;
wire v_EXEC2_3170_out0;
wire v_EXEC2_3171_out0;
wire v_EXEC2_3241_out0;
wire v_EXEC2_3242_out0;
wire v_EXEC2_441_out0;
wire v_EXEC2_442_out0;
wire v_EXEC2_7181_out0;
wire v_EXEC2_7182_out0;
wire v_EXP1_13488_out0;
wire v_EXP1_13489_out0;
wire v_FLAOTING_INSTRUCTION_1859_out0;
wire v_FLAOTING_INSTRUCTION_1860_out0;
wire v_FLOATING_EN_ALU_634_out0;
wire v_FLOATING_EN_ALU_635_out0;
wire v_FLOATING_INSTRUCTION_10391_out0;
wire v_FLOATING_INSTRUCTION_10392_out0;
wire v_FLOATING_INS_13797_out0;
wire v_FLOATING_INS_13798_out0;
wire v_FLOAT_4603_out0;
wire v_FLOAT_4604_out0;
wire v_FLOAT_7676_out0;
wire v_FLOAT_7677_out0;
wire v_FLOAT_INST16_13443_out0;
wire v_FLOAT_INST16_13444_out0;
wire v_FLOAT_INST_2955_out0;
wire v_FLOAT_INST_2956_out0;
wire v_G10_10694_out0;
wire v_G10_10711_out0;
wire v_G10_130_out0;
wire v_G10_131_out0;
wire v_G10_13215_out0;
wire v_G10_13216_out0;
wire v_G10_13217_out0;
wire v_G10_13218_out0;
wire v_G10_1755_out0;
wire v_G10_1756_out0;
wire v_G10_1943_out0;
wire v_G10_1944_out0;
wire v_G10_1945_out0;
wire v_G10_1946_out0;
wire v_G10_2632_out0;
wire v_G10_2633_out0;
wire v_G10_2640_out0;
wire v_G10_2641_out0;
wire v_G10_2642_out0;
wire v_G10_2643_out0;
wire v_G10_4479_out0;
wire v_G10_4480_out0;
wire v_G10_602_out0;
wire v_G10_6975_out0;
wire v_G10_6976_out0;
wire v_G10_6977_out0;
wire v_G10_6978_out0;
wire v_G10_6979_out0;
wire v_G10_6980_out0;
wire v_G10_6981_out0;
wire v_G10_6982_out0;
wire v_G10_6983_out0;
wire v_G10_6984_out0;
wire v_G10_6985_out0;
wire v_G10_6986_out0;
wire v_G10_6987_out0;
wire v_G10_6988_out0;
wire v_G10_6989_out0;
wire v_G10_6990_out0;
wire v_G10_6991_out0;
wire v_G10_6992_out0;
wire v_G10_6993_out0;
wire v_G10_6994_out0;
wire v_G10_6995_out0;
wire v_G10_6996_out0;
wire v_G10_6997_out0;
wire v_G10_6998_out0;
wire v_G10_6999_out0;
wire v_G10_7000_out0;
wire v_G10_7001_out0;
wire v_G10_7002_out0;
wire v_G10_7003_out0;
wire v_G10_7004_out0;
wire v_G11_11165_out0;
wire v_G11_11166_out0;
wire v_G11_13342_out0;
wire v_G11_13343_out0;
wire v_G11_13344_out0;
wire v_G11_13345_out0;
wire v_G11_13439_out0;
wire v_G11_13440_out0;
wire v_G11_2550_out0;
wire v_G11_2551_out0;
wire v_G11_2626_out0;
wire v_G11_2627_out0;
wire v_G11_2937_out0;
wire v_G11_2938_out0;
wire v_G11_2939_out0;
wire v_G11_2940_out0;
wire v_G11_651_out0;
wire v_G11_652_out0;
wire v_G11_653_out0;
wire v_G11_654_out0;
wire v_G11_655_out0;
wire v_G11_656_out0;
wire v_G11_657_out0;
wire v_G11_658_out0;
wire v_G11_659_out0;
wire v_G11_660_out0;
wire v_G11_661_out0;
wire v_G11_662_out0;
wire v_G11_663_out0;
wire v_G11_664_out0;
wire v_G11_665_out0;
wire v_G11_666_out0;
wire v_G11_667_out0;
wire v_G11_668_out0;
wire v_G11_669_out0;
wire v_G11_670_out0;
wire v_G11_671_out0;
wire v_G11_672_out0;
wire v_G11_673_out0;
wire v_G11_674_out0;
wire v_G11_675_out0;
wire v_G11_676_out0;
wire v_G11_677_out0;
wire v_G11_678_out0;
wire v_G11_679_out0;
wire v_G11_680_out0;
wire v_G11_8652_out0;
wire v_G12_10321_out0;
wire v_G12_10322_out0;
wire v_G12_10688_out0;
wire v_G12_10689_out0;
wire v_G12_10690_out0;
wire v_G12_10691_out0;
wire v_G12_13221_out0;
wire v_G12_13222_out0;
wire v_G12_13223_out0;
wire v_G12_13224_out0;
wire v_G12_13225_out0;
wire v_G12_13226_out0;
wire v_G12_13227_out0;
wire v_G12_13228_out0;
wire v_G12_13229_out0;
wire v_G12_13230_out0;
wire v_G12_13231_out0;
wire v_G12_13232_out0;
wire v_G12_13233_out0;
wire v_G12_13234_out0;
wire v_G12_13235_out0;
wire v_G12_13236_out0;
wire v_G12_13237_out0;
wire v_G12_13238_out0;
wire v_G12_13239_out0;
wire v_G12_13240_out0;
wire v_G12_13241_out0;
wire v_G12_13242_out0;
wire v_G12_13243_out0;
wire v_G12_13244_out0;
wire v_G12_13245_out0;
wire v_G12_13246_out0;
wire v_G12_13247_out0;
wire v_G12_13248_out0;
wire v_G12_13249_out0;
wire v_G12_13250_out0;
wire v_G12_2270_out0;
wire v_G12_3345_out0;
wire v_G12_3346_out0;
wire v_G12_3347_out0;
wire v_G12_3348_out0;
wire v_G12_4699_out0;
wire v_G12_4700_out0;
wire v_G13_13352_out0;
wire v_G13_13353_out0;
wire v_G13_13354_out0;
wire v_G13_13355_out0;
wire v_G13_13356_out0;
wire v_G13_13357_out0;
wire v_G13_13358_out0;
wire v_G13_13359_out0;
wire v_G13_13360_out0;
wire v_G13_13361_out0;
wire v_G13_13362_out0;
wire v_G13_13363_out0;
wire v_G13_13364_out0;
wire v_G13_13365_out0;
wire v_G13_13366_out0;
wire v_G13_13367_out0;
wire v_G13_13368_out0;
wire v_G13_13369_out0;
wire v_G13_13370_out0;
wire v_G13_13371_out0;
wire v_G13_13372_out0;
wire v_G13_13373_out0;
wire v_G13_13374_out0;
wire v_G13_13375_out0;
wire v_G13_13376_out0;
wire v_G13_13377_out0;
wire v_G13_13378_out0;
wire v_G13_13379_out0;
wire v_G13_13380_out0;
wire v_G13_13381_out0;
wire v_G13_4705_out0;
wire v_G13_4706_out0;
wire v_G13_4707_out0;
wire v_G13_4708_out0;
wire v_G13_642_out0;
wire v_G13_643_out0;
wire v_G13_644_out0;
wire v_G13_645_out0;
wire v_G13_7083_out0;
wire v_G13_7084_out0;
wire v_G14_10407_out0;
wire v_G14_10408_out0;
wire v_G14_1178_out0;
wire v_G14_1179_out0;
wire v_G14_13268_out0;
wire v_G14_13269_out0;
wire v_G14_13672_out0;
wire v_G14_13673_out0;
wire v_G14_13674_out0;
wire v_G14_13675_out0;
wire v_G14_13676_out0;
wire v_G14_13677_out0;
wire v_G14_13678_out0;
wire v_G14_13679_out0;
wire v_G14_13680_out0;
wire v_G14_13681_out0;
wire v_G14_13682_out0;
wire v_G14_13683_out0;
wire v_G14_13684_out0;
wire v_G14_13685_out0;
wire v_G14_13686_out0;
wire v_G14_13687_out0;
wire v_G14_13688_out0;
wire v_G14_13689_out0;
wire v_G14_13690_out0;
wire v_G14_13691_out0;
wire v_G14_13692_out0;
wire v_G14_13693_out0;
wire v_G14_13694_out0;
wire v_G14_13695_out0;
wire v_G14_13696_out0;
wire v_G14_13697_out0;
wire v_G14_13698_out0;
wire v_G14_13699_out0;
wire v_G14_13700_out0;
wire v_G14_13701_out0;
wire v_G14_4533_out0;
wire v_G14_4534_out0;
wire v_G14_4535_out0;
wire v_G14_4536_out0;
wire v_G14_615_out0;
wire v_G14_616_out0;
wire v_G14_617_out0;
wire v_G14_618_out0;
wire v_G15_132_out0;
wire v_G15_133_out0;
wire v_G15_134_out0;
wire v_G15_135_out0;
wire v_G15_136_out0;
wire v_G15_137_out0;
wire v_G15_138_out0;
wire v_G15_139_out0;
wire v_G15_140_out0;
wire v_G15_141_out0;
wire v_G15_142_out0;
wire v_G15_143_out0;
wire v_G15_144_out0;
wire v_G15_145_out0;
wire v_G15_146_out0;
wire v_G15_147_out0;
wire v_G15_148_out0;
wire v_G15_149_out0;
wire v_G15_150_out0;
wire v_G15_151_out0;
wire v_G15_152_out0;
wire v_G15_153_out0;
wire v_G15_154_out0;
wire v_G15_155_out0;
wire v_G15_156_out0;
wire v_G15_157_out0;
wire v_G15_158_out0;
wire v_G15_159_out0;
wire v_G15_160_out0;
wire v_G15_161_out0;
wire v_G15_1814_out0;
wire v_G15_1815_out0;
wire v_G15_1816_out0;
wire v_G15_1817_out0;
wire v_G15_1855_out0;
wire v_G15_1856_out0;
wire v_G15_4654_out0;
wire v_G15_4655_out0;
wire v_G15_4656_out0;
wire v_G15_4657_out0;
wire v_G16_10906_out0;
wire v_G16_10907_out0;
wire v_G16_10908_out0;
wire v_G16_10909_out0;
wire v_G16_11034_out0;
wire v_G16_11035_out0;
wire v_G16_11036_out0;
wire v_G16_11037_out0;
wire v_G16_13183_out0;
wire v_G16_13184_out0;
wire v_G16_13185_out0;
wire v_G16_13186_out0;
wire v_G16_13187_out0;
wire v_G16_13188_out0;
wire v_G16_13189_out0;
wire v_G16_13190_out0;
wire v_G16_13191_out0;
wire v_G16_13192_out0;
wire v_G16_13193_out0;
wire v_G16_13194_out0;
wire v_G16_13195_out0;
wire v_G16_13196_out0;
wire v_G16_13197_out0;
wire v_G16_13198_out0;
wire v_G16_13199_out0;
wire v_G16_13200_out0;
wire v_G16_13201_out0;
wire v_G16_13202_out0;
wire v_G16_13203_out0;
wire v_G16_13204_out0;
wire v_G16_13205_out0;
wire v_G16_13206_out0;
wire v_G16_13207_out0;
wire v_G16_13208_out0;
wire v_G16_13209_out0;
wire v_G16_13210_out0;
wire v_G16_13211_out0;
wire v_G16_13212_out0;
wire v_G16_13388_out0;
wire v_G16_13389_out0;
wire v_G16_2310_out0;
wire v_G16_2311_out0;
wire v_G16_3024_out0;
wire v_G16_7701_out0;
wire v_G17_10710_out0;
wire v_G17_1903_out0;
wire v_G18_10489_out0;
wire v_G18_11204_out0;
wire v_G18_11205_out0;
wire v_G18_2407_out0;
wire v_G18_2408_out0;
wire v_G18_567_out0;
wire v_G18_8799_out0;
wire v_G18_8800_out0;
wire v_G18_8801_out0;
wire v_G18_8802_out0;
wire v_G19_10327_out0;
wire v_G19_10328_out0;
wire v_G19_3860_out0;
wire v_G19_4663_out0;
wire v_G19_4664_out0;
wire v_G1_10476_out0;
wire v_G1_10477_out0;
wire v_G1_10478_out0;
wire v_G1_10757_out0;
wire v_G1_10758_out0;
wire v_G1_10810_out0;
wire v_G1_11157_out0;
wire v_G1_11158_out0;
wire v_G1_1167_out0;
wire v_G1_1168_out0;
wire v_G1_1191_out0;
wire v_G1_1192_out0;
wire v_G1_13757_out0;
wire v_G1_13758_out0;
wire v_G1_13759_out0;
wire v_G1_13760_out0;
wire v_G1_13776_out0;
wire v_G1_13777_out0;
wire v_G1_1879_out0;
wire v_G1_1880_out0;
wire v_G1_1881_out0;
wire v_G1_1882_out0;
wire v_G1_1909_out0;
wire v_G1_1910_out0;
wire v_G1_1911_out0;
wire v_G1_1912_out0;
wire v_G1_1913_out0;
wire v_G1_1914_out0;
wire v_G1_1915_out0;
wire v_G1_1916_out0;
wire v_G1_1917_out0;
wire v_G1_1918_out0;
wire v_G1_1919_out0;
wire v_G1_1920_out0;
wire v_G1_1921_out0;
wire v_G1_1922_out0;
wire v_G1_1923_out0;
wire v_G1_1924_out0;
wire v_G1_1925_out0;
wire v_G1_1926_out0;
wire v_G1_1927_out0;
wire v_G1_1928_out0;
wire v_G1_1929_out0;
wire v_G1_1930_out0;
wire v_G1_1931_out0;
wire v_G1_1932_out0;
wire v_G1_1933_out0;
wire v_G1_1934_out0;
wire v_G1_1935_out0;
wire v_G1_1936_out0;
wire v_G1_1937_out0;
wire v_G1_1938_out0;
wire v_G1_2225_out0;
wire v_G1_2226_out0;
wire v_G1_2354_out0;
wire v_G1_2700_out0;
wire v_G1_2701_out0;
wire v_G1_2702_out0;
wire v_G1_2703_out0;
wire v_G1_2704_out0;
wire v_G1_2705_out0;
wire v_G1_2706_out0;
wire v_G1_2707_out0;
wire v_G1_2708_out0;
wire v_G1_2709_out0;
wire v_G1_2710_out0;
wire v_G1_2711_out0;
wire v_G1_2712_out0;
wire v_G1_2713_out0;
wire v_G1_2714_out0;
wire v_G1_2715_out0;
wire v_G1_277_out0;
wire v_G1_289_out0;
wire v_G1_290_out0;
wire v_G1_2911_out0;
wire v_G1_3018_out0;
wire v_G1_3019_out0;
wire v_G1_3995_out0;
wire v_G1_3996_out0;
wire v_G1_3997_out0;
wire v_G1_3998_out0;
wire v_G1_3999_out0;
wire v_G1_4000_out0;
wire v_G1_4001_out0;
wire v_G1_4002_out0;
wire v_G1_4003_out0;
wire v_G1_4004_out0;
wire v_G1_4005_out0;
wire v_G1_4006_out0;
wire v_G1_4007_out0;
wire v_G1_4008_out0;
wire v_G1_4009_out0;
wire v_G1_4010_out0;
wire v_G1_4011_out0;
wire v_G1_4012_out0;
wire v_G1_4013_out0;
wire v_G1_4014_out0;
wire v_G1_4015_out0;
wire v_G1_4016_out0;
wire v_G1_4017_out0;
wire v_G1_4018_out0;
wire v_G1_4019_out0;
wire v_G1_4020_out0;
wire v_G1_4021_out0;
wire v_G1_4022_out0;
wire v_G1_4023_out0;
wire v_G1_4024_out0;
wire v_G1_4025_out0;
wire v_G1_4026_out0;
wire v_G1_4027_out0;
wire v_G1_4028_out0;
wire v_G1_4029_out0;
wire v_G1_4030_out0;
wire v_G1_4031_out0;
wire v_G1_4032_out0;
wire v_G1_4033_out0;
wire v_G1_4034_out0;
wire v_G1_4035_out0;
wire v_G1_4036_out0;
wire v_G1_4037_out0;
wire v_G1_4038_out0;
wire v_G1_4039_out0;
wire v_G1_4040_out0;
wire v_G1_4041_out0;
wire v_G1_4042_out0;
wire v_G1_4043_out0;
wire v_G1_4044_out0;
wire v_G1_4045_out0;
wire v_G1_4046_out0;
wire v_G1_4047_out0;
wire v_G1_4048_out0;
wire v_G1_4049_out0;
wire v_G1_4050_out0;
wire v_G1_4051_out0;
wire v_G1_4052_out0;
wire v_G1_4053_out0;
wire v_G1_4054_out0;
wire v_G1_4055_out0;
wire v_G1_4056_out0;
wire v_G1_4057_out0;
wire v_G1_4058_out0;
wire v_G1_4059_out0;
wire v_G1_4060_out0;
wire v_G1_4061_out0;
wire v_G1_4062_out0;
wire v_G1_4063_out0;
wire v_G1_4064_out0;
wire v_G1_4065_out0;
wire v_G1_4066_out0;
wire v_G1_4067_out0;
wire v_G1_4068_out0;
wire v_G1_4069_out0;
wire v_G1_4070_out0;
wire v_G1_4071_out0;
wire v_G1_4072_out0;
wire v_G1_4073_out0;
wire v_G1_4074_out0;
wire v_G1_4075_out0;
wire v_G1_4076_out0;
wire v_G1_4077_out0;
wire v_G1_4078_out0;
wire v_G1_4079_out0;
wire v_G1_4080_out0;
wire v_G1_4081_out0;
wire v_G1_4082_out0;
wire v_G1_4083_out0;
wire v_G1_4084_out0;
wire v_G1_4085_out0;
wire v_G1_4086_out0;
wire v_G1_4087_out0;
wire v_G1_4088_out0;
wire v_G1_4089_out0;
wire v_G1_4090_out0;
wire v_G1_4091_out0;
wire v_G1_4092_out0;
wire v_G1_4093_out0;
wire v_G1_4094_out0;
wire v_G1_4095_out0;
wire v_G1_4096_out0;
wire v_G1_4097_out0;
wire v_G1_4098_out0;
wire v_G1_4099_out0;
wire v_G1_4100_out0;
wire v_G1_4101_out0;
wire v_G1_4102_out0;
wire v_G1_4103_out0;
wire v_G1_4104_out0;
wire v_G1_4105_out0;
wire v_G1_4106_out0;
wire v_G1_4107_out0;
wire v_G1_4108_out0;
wire v_G1_4109_out0;
wire v_G1_4110_out0;
wire v_G1_4111_out0;
wire v_G1_4112_out0;
wire v_G1_4113_out0;
wire v_G1_4114_out0;
wire v_G1_4115_out0;
wire v_G1_4116_out0;
wire v_G1_4117_out0;
wire v_G1_4118_out0;
wire v_G1_4119_out0;
wire v_G1_4120_out0;
wire v_G1_4121_out0;
wire v_G1_4122_out0;
wire v_G1_4123_out0;
wire v_G1_4124_out0;
wire v_G1_4125_out0;
wire v_G1_4126_out0;
wire v_G1_4127_out0;
wire v_G1_4128_out0;
wire v_G1_4129_out0;
wire v_G1_4130_out0;
wire v_G1_4131_out0;
wire v_G1_4132_out0;
wire v_G1_4133_out0;
wire v_G1_4134_out0;
wire v_G1_4135_out0;
wire v_G1_4136_out0;
wire v_G1_4137_out0;
wire v_G1_4138_out0;
wire v_G1_4139_out0;
wire v_G1_4140_out0;
wire v_G1_4141_out0;
wire v_G1_4142_out0;
wire v_G1_4143_out0;
wire v_G1_4144_out0;
wire v_G1_4145_out0;
wire v_G1_4146_out0;
wire v_G1_4147_out0;
wire v_G1_4148_out0;
wire v_G1_4149_out0;
wire v_G1_4150_out0;
wire v_G1_4151_out0;
wire v_G1_4152_out0;
wire v_G1_4153_out0;
wire v_G1_4154_out0;
wire v_G1_4155_out0;
wire v_G1_4156_out0;
wire v_G1_4157_out0;
wire v_G1_4158_out0;
wire v_G1_4159_out0;
wire v_G1_4160_out0;
wire v_G1_4161_out0;
wire v_G1_4162_out0;
wire v_G1_4163_out0;
wire v_G1_4164_out0;
wire v_G1_4165_out0;
wire v_G1_4166_out0;
wire v_G1_4167_out0;
wire v_G1_4168_out0;
wire v_G1_4169_out0;
wire v_G1_4170_out0;
wire v_G1_4171_out0;
wire v_G1_4172_out0;
wire v_G1_4173_out0;
wire v_G1_4174_out0;
wire v_G1_4175_out0;
wire v_G1_4176_out0;
wire v_G1_4177_out0;
wire v_G1_4178_out0;
wire v_G1_4179_out0;
wire v_G1_4180_out0;
wire v_G1_4181_out0;
wire v_G1_4182_out0;
wire v_G1_4183_out0;
wire v_G1_4184_out0;
wire v_G1_4185_out0;
wire v_G1_4186_out0;
wire v_G1_4187_out0;
wire v_G1_4188_out0;
wire v_G1_4189_out0;
wire v_G1_4190_out0;
wire v_G1_4191_out0;
wire v_G1_4192_out0;
wire v_G1_4193_out0;
wire v_G1_4194_out0;
wire v_G1_4195_out0;
wire v_G1_4196_out0;
wire v_G1_4197_out0;
wire v_G1_4198_out0;
wire v_G1_4199_out0;
wire v_G1_4200_out0;
wire v_G1_4201_out0;
wire v_G1_4202_out0;
wire v_G1_4203_out0;
wire v_G1_4204_out0;
wire v_G1_4205_out0;
wire v_G1_4206_out0;
wire v_G1_4207_out0;
wire v_G1_4208_out0;
wire v_G1_4209_out0;
wire v_G1_4210_out0;
wire v_G1_4211_out0;
wire v_G1_4212_out0;
wire v_G1_4213_out0;
wire v_G1_4214_out0;
wire v_G1_4215_out0;
wire v_G1_4216_out0;
wire v_G1_4217_out0;
wire v_G1_4218_out0;
wire v_G1_4219_out0;
wire v_G1_4220_out0;
wire v_G1_4221_out0;
wire v_G1_4222_out0;
wire v_G1_4223_out0;
wire v_G1_4224_out0;
wire v_G1_4225_out0;
wire v_G1_4226_out0;
wire v_G1_4227_out0;
wire v_G1_4228_out0;
wire v_G1_4229_out0;
wire v_G1_4230_out0;
wire v_G1_4231_out0;
wire v_G1_4232_out0;
wire v_G1_4233_out0;
wire v_G1_4234_out0;
wire v_G1_4235_out0;
wire v_G1_4236_out0;
wire v_G1_4237_out0;
wire v_G1_4238_out0;
wire v_G1_4239_out0;
wire v_G1_4240_out0;
wire v_G1_4241_out0;
wire v_G1_4242_out0;
wire v_G1_4243_out0;
wire v_G1_4244_out0;
wire v_G1_4245_out0;
wire v_G1_4246_out0;
wire v_G1_4247_out0;
wire v_G1_4248_out0;
wire v_G1_4249_out0;
wire v_G1_4250_out0;
wire v_G1_4251_out0;
wire v_G1_4252_out0;
wire v_G1_4253_out0;
wire v_G1_4254_out0;
wire v_G1_4255_out0;
wire v_G1_4256_out0;
wire v_G1_4257_out0;
wire v_G1_4258_out0;
wire v_G1_4259_out0;
wire v_G1_4260_out0;
wire v_G1_4261_out0;
wire v_G1_4262_out0;
wire v_G1_4263_out0;
wire v_G1_4264_out0;
wire v_G1_4265_out0;
wire v_G1_4266_out0;
wire v_G1_4267_out0;
wire v_G1_4268_out0;
wire v_G1_4269_out0;
wire v_G1_4270_out0;
wire v_G1_4271_out0;
wire v_G1_4272_out0;
wire v_G1_4273_out0;
wire v_G1_4274_out0;
wire v_G1_4275_out0;
wire v_G1_4276_out0;
wire v_G1_4277_out0;
wire v_G1_4278_out0;
wire v_G1_4279_out0;
wire v_G1_4280_out0;
wire v_G1_4281_out0;
wire v_G1_4282_out0;
wire v_G1_4283_out0;
wire v_G1_4284_out0;
wire v_G1_4285_out0;
wire v_G1_4286_out0;
wire v_G1_4287_out0;
wire v_G1_4288_out0;
wire v_G1_4289_out0;
wire v_G1_4290_out0;
wire v_G1_4291_out0;
wire v_G1_4292_out0;
wire v_G1_4293_out0;
wire v_G1_4294_out0;
wire v_G1_4295_out0;
wire v_G1_4296_out0;
wire v_G1_4297_out0;
wire v_G1_4298_out0;
wire v_G1_4299_out0;
wire v_G1_4300_out0;
wire v_G1_4301_out0;
wire v_G1_4302_out0;
wire v_G1_4303_out0;
wire v_G1_4304_out0;
wire v_G1_4305_out0;
wire v_G1_4306_out0;
wire v_G1_4307_out0;
wire v_G1_4308_out0;
wire v_G1_4309_out0;
wire v_G1_4310_out0;
wire v_G1_4311_out0;
wire v_G1_4312_out0;
wire v_G1_4313_out0;
wire v_G1_4314_out0;
wire v_G1_4315_out0;
wire v_G1_4316_out0;
wire v_G1_4317_out0;
wire v_G1_4318_out0;
wire v_G1_4319_out0;
wire v_G1_4320_out0;
wire v_G1_4321_out0;
wire v_G1_4322_out0;
wire v_G1_4323_out0;
wire v_G1_4324_out0;
wire v_G1_4325_out0;
wire v_G1_4326_out0;
wire v_G1_4327_out0;
wire v_G1_4328_out0;
wire v_G1_4329_out0;
wire v_G1_4330_out0;
wire v_G1_4331_out0;
wire v_G1_4332_out0;
wire v_G1_4333_out0;
wire v_G1_4334_out0;
wire v_G1_4335_out0;
wire v_G1_4336_out0;
wire v_G1_4337_out0;
wire v_G1_4338_out0;
wire v_G1_4339_out0;
wire v_G1_4340_out0;
wire v_G1_4341_out0;
wire v_G1_4342_out0;
wire v_G1_4343_out0;
wire v_G1_4344_out0;
wire v_G1_4345_out0;
wire v_G1_4346_out0;
wire v_G1_4347_out0;
wire v_G1_4348_out0;
wire v_G1_4349_out0;
wire v_G1_4350_out0;
wire v_G1_4351_out0;
wire v_G1_4352_out0;
wire v_G1_4353_out0;
wire v_G1_4354_out0;
wire v_G1_4355_out0;
wire v_G1_4356_out0;
wire v_G1_4357_out0;
wire v_G1_4358_out0;
wire v_G1_4359_out0;
wire v_G1_4360_out0;
wire v_G1_4361_out0;
wire v_G1_4362_out0;
wire v_G1_4363_out0;
wire v_G1_4364_out0;
wire v_G1_4365_out0;
wire v_G1_4366_out0;
wire v_G1_4367_out0;
wire v_G1_4368_out0;
wire v_G1_4369_out0;
wire v_G1_4370_out0;
wire v_G1_4371_out0;
wire v_G1_4372_out0;
wire v_G1_4373_out0;
wire v_G1_4374_out0;
wire v_G1_4375_out0;
wire v_G1_4376_out0;
wire v_G1_4377_out0;
wire v_G1_4378_out0;
wire v_G1_4379_out0;
wire v_G1_4380_out0;
wire v_G1_4381_out0;
wire v_G1_4382_out0;
wire v_G1_4383_out0;
wire v_G1_4384_out0;
wire v_G1_4385_out0;
wire v_G1_4386_out0;
wire v_G1_4387_out0;
wire v_G1_4388_out0;
wire v_G1_4389_out0;
wire v_G1_4390_out0;
wire v_G1_4391_out0;
wire v_G1_4392_out0;
wire v_G1_4393_out0;
wire v_G1_4394_out0;
wire v_G1_4395_out0;
wire v_G1_4396_out0;
wire v_G1_4397_out0;
wire v_G1_4398_out0;
wire v_G1_4399_out0;
wire v_G1_4400_out0;
wire v_G1_4401_out0;
wire v_G1_4402_out0;
wire v_G1_4403_out0;
wire v_G1_4404_out0;
wire v_G1_4405_out0;
wire v_G1_4406_out0;
wire v_G1_4407_out0;
wire v_G1_4408_out0;
wire v_G1_4409_out0;
wire v_G1_4410_out0;
wire v_G1_4411_out0;
wire v_G1_4412_out0;
wire v_G1_4413_out0;
wire v_G1_4414_out0;
wire v_G1_4415_out0;
wire v_G1_4416_out0;
wire v_G1_4417_out0;
wire v_G1_4418_out0;
wire v_G1_4419_out0;
wire v_G1_4420_out0;
wire v_G1_4421_out0;
wire v_G1_4422_out0;
wire v_G1_4423_out0;
wire v_G1_4424_out0;
wire v_G1_4425_out0;
wire v_G1_4426_out0;
wire v_G1_4427_out0;
wire v_G1_4428_out0;
wire v_G1_4429_out0;
wire v_G1_4430_out0;
wire v_G1_4431_out0;
wire v_G1_4432_out0;
wire v_G1_4433_out0;
wire v_G1_4434_out0;
wire v_G1_4435_out0;
wire v_G1_4436_out0;
wire v_G1_4437_out0;
wire v_G1_4438_out0;
wire v_G1_4439_out0;
wire v_G1_4440_out0;
wire v_G1_4441_out0;
wire v_G1_4442_out0;
wire v_G1_646_out0;
wire v_G1_647_out0;
wire v_G1_7717_out0;
wire v_G1_7718_out0;
wire v_G1_7719_out0;
wire v_G1_7720_out0;
wire v_G1_7721_out0;
wire v_G1_7722_out0;
wire v_G1_7723_out0;
wire v_G1_7724_out0;
wire v_G1_7725_out0;
wire v_G1_7726_out0;
wire v_G1_7727_out0;
wire v_G1_7728_out0;
wire v_G1_7729_out0;
wire v_G1_7730_out0;
wire v_G1_7731_out0;
wire v_G1_7732_out0;
wire v_G1_7733_out0;
wire v_G1_7734_out0;
wire v_G1_7735_out0;
wire v_G1_7736_out0;
wire v_G1_7737_out0;
wire v_G1_7738_out0;
wire v_G1_7739_out0;
wire v_G1_7740_out0;
wire v_G1_7741_out0;
wire v_G1_7742_out0;
wire v_G1_7743_out0;
wire v_G1_7744_out0;
wire v_G1_7745_out0;
wire v_G1_7746_out0;
wire v_G1_7747_out0;
wire v_G1_7748_out0;
wire v_G1_7749_out0;
wire v_G1_7750_out0;
wire v_G1_7751_out0;
wire v_G1_7752_out0;
wire v_G1_7753_out0;
wire v_G1_7754_out0;
wire v_G1_7755_out0;
wire v_G1_7756_out0;
wire v_G1_7757_out0;
wire v_G1_7758_out0;
wire v_G1_7759_out0;
wire v_G1_7760_out0;
wire v_G1_7761_out0;
wire v_G1_7762_out0;
wire v_G1_7763_out0;
wire v_G1_7764_out0;
wire v_G1_7765_out0;
wire v_G1_7766_out0;
wire v_G1_7767_out0;
wire v_G1_7768_out0;
wire v_G1_7769_out0;
wire v_G1_7770_out0;
wire v_G1_7771_out0;
wire v_G1_7772_out0;
wire v_G1_7773_out0;
wire v_G1_7774_out0;
wire v_G1_7775_out0;
wire v_G1_7776_out0;
wire v_G1_7777_out0;
wire v_G1_7778_out0;
wire v_G1_7779_out0;
wire v_G1_7780_out0;
wire v_G1_7781_out0;
wire v_G1_7782_out0;
wire v_G1_7783_out0;
wire v_G1_7784_out0;
wire v_G1_7785_out0;
wire v_G1_7786_out0;
wire v_G1_7787_out0;
wire v_G1_7788_out0;
wire v_G1_7789_out0;
wire v_G1_7790_out0;
wire v_G1_7791_out0;
wire v_G1_7792_out0;
wire v_G1_7793_out0;
wire v_G1_7794_out0;
wire v_G1_7795_out0;
wire v_G1_7796_out0;
wire v_G1_7797_out0;
wire v_G1_7798_out0;
wire v_G1_7799_out0;
wire v_G1_7800_out0;
wire v_G1_7801_out0;
wire v_G1_7802_out0;
wire v_G1_7803_out0;
wire v_G1_7804_out0;
wire v_G1_7805_out0;
wire v_G1_7806_out0;
wire v_G1_7807_out0;
wire v_G1_7808_out0;
wire v_G1_7809_out0;
wire v_G1_7810_out0;
wire v_G1_7811_out0;
wire v_G1_7812_out0;
wire v_G1_7813_out0;
wire v_G1_7814_out0;
wire v_G1_7815_out0;
wire v_G1_7816_out0;
wire v_G1_7817_out0;
wire v_G1_7818_out0;
wire v_G1_7819_out0;
wire v_G1_7820_out0;
wire v_G1_7821_out0;
wire v_G1_7822_out0;
wire v_G1_7823_out0;
wire v_G1_7824_out0;
wire v_G1_7825_out0;
wire v_G1_7826_out0;
wire v_G1_7827_out0;
wire v_G1_7828_out0;
wire v_G1_7829_out0;
wire v_G1_7830_out0;
wire v_G1_7831_out0;
wire v_G1_7832_out0;
wire v_G1_7833_out0;
wire v_G1_7834_out0;
wire v_G1_7835_out0;
wire v_G1_7836_out0;
wire v_G1_7837_out0;
wire v_G1_7838_out0;
wire v_G1_7839_out0;
wire v_G1_7840_out0;
wire v_G1_7841_out0;
wire v_G1_7842_out0;
wire v_G1_7843_out0;
wire v_G1_7844_out0;
wire v_G1_7845_out0;
wire v_G1_7846_out0;
wire v_G1_7847_out0;
wire v_G1_7848_out0;
wire v_G1_7849_out0;
wire v_G1_7850_out0;
wire v_G1_7851_out0;
wire v_G1_7852_out0;
wire v_G1_7853_out0;
wire v_G1_7854_out0;
wire v_G1_7855_out0;
wire v_G1_7856_out0;
wire v_G1_7857_out0;
wire v_G1_7858_out0;
wire v_G1_7859_out0;
wire v_G1_7860_out0;
wire v_G1_7861_out0;
wire v_G1_7862_out0;
wire v_G1_7863_out0;
wire v_G1_7864_out0;
wire v_G1_7865_out0;
wire v_G1_7866_out0;
wire v_G1_7867_out0;
wire v_G1_7868_out0;
wire v_G1_7869_out0;
wire v_G1_7870_out0;
wire v_G1_7871_out0;
wire v_G1_7872_out0;
wire v_G1_7873_out0;
wire v_G1_7874_out0;
wire v_G1_7875_out0;
wire v_G1_7876_out0;
wire v_G1_7877_out0;
wire v_G1_7878_out0;
wire v_G1_7879_out0;
wire v_G1_7880_out0;
wire v_G1_7881_out0;
wire v_G1_7882_out0;
wire v_G1_7883_out0;
wire v_G1_7884_out0;
wire v_G1_7885_out0;
wire v_G1_7886_out0;
wire v_G1_7887_out0;
wire v_G1_7888_out0;
wire v_G1_7889_out0;
wire v_G1_7890_out0;
wire v_G1_7891_out0;
wire v_G1_7892_out0;
wire v_G1_7893_out0;
wire v_G1_7894_out0;
wire v_G1_7895_out0;
wire v_G1_7896_out0;
wire v_G1_7897_out0;
wire v_G1_7898_out0;
wire v_G1_7899_out0;
wire v_G1_7900_out0;
wire v_G1_7901_out0;
wire v_G1_7902_out0;
wire v_G1_7903_out0;
wire v_G1_7904_out0;
wire v_G1_7905_out0;
wire v_G1_7906_out0;
wire v_G1_7907_out0;
wire v_G1_7908_out0;
wire v_G1_7909_out0;
wire v_G1_7910_out0;
wire v_G1_7911_out0;
wire v_G1_7912_out0;
wire v_G1_7913_out0;
wire v_G1_7914_out0;
wire v_G1_7915_out0;
wire v_G1_7916_out0;
wire v_G1_7917_out0;
wire v_G1_7918_out0;
wire v_G1_7919_out0;
wire v_G1_7920_out0;
wire v_G1_7921_out0;
wire v_G1_7922_out0;
wire v_G1_7923_out0;
wire v_G1_7924_out0;
wire v_G1_7925_out0;
wire v_G1_7926_out0;
wire v_G1_7927_out0;
wire v_G1_7928_out0;
wire v_G1_7929_out0;
wire v_G1_7930_out0;
wire v_G1_7931_out0;
wire v_G1_7932_out0;
wire v_G1_7933_out0;
wire v_G1_7934_out0;
wire v_G1_7935_out0;
wire v_G1_7936_out0;
wire v_G1_7937_out0;
wire v_G1_7938_out0;
wire v_G1_7939_out0;
wire v_G1_7940_out0;
wire v_G1_7941_out0;
wire v_G1_7942_out0;
wire v_G1_7943_out0;
wire v_G1_7944_out0;
wire v_G1_7945_out0;
wire v_G1_7946_out0;
wire v_G1_7947_out0;
wire v_G1_7948_out0;
wire v_G1_7949_out0;
wire v_G1_7950_out0;
wire v_G1_7951_out0;
wire v_G1_7952_out0;
wire v_G1_7953_out0;
wire v_G1_7954_out0;
wire v_G1_7955_out0;
wire v_G1_7956_out0;
wire v_G1_7957_out0;
wire v_G1_7958_out0;
wire v_G1_7959_out0;
wire v_G1_7960_out0;
wire v_G1_7961_out0;
wire v_G1_7962_out0;
wire v_G1_7963_out0;
wire v_G1_7964_out0;
wire v_G1_7965_out0;
wire v_G1_7966_out0;
wire v_G1_7967_out0;
wire v_G1_7968_out0;
wire v_G1_7969_out0;
wire v_G1_7970_out0;
wire v_G1_7971_out0;
wire v_G1_7972_out0;
wire v_G1_7973_out0;
wire v_G1_7974_out0;
wire v_G1_7975_out0;
wire v_G1_7976_out0;
wire v_G1_7977_out0;
wire v_G1_7978_out0;
wire v_G1_7979_out0;
wire v_G1_7980_out0;
wire v_G1_7981_out0;
wire v_G1_7982_out0;
wire v_G1_7983_out0;
wire v_G1_7984_out0;
wire v_G1_7985_out0;
wire v_G1_7986_out0;
wire v_G1_7987_out0;
wire v_G1_7988_out0;
wire v_G1_7989_out0;
wire v_G1_7990_out0;
wire v_G1_7991_out0;
wire v_G1_7992_out0;
wire v_G1_7993_out0;
wire v_G1_7994_out0;
wire v_G1_7995_out0;
wire v_G1_7996_out0;
wire v_G1_7997_out0;
wire v_G1_7998_out0;
wire v_G1_7999_out0;
wire v_G1_8000_out0;
wire v_G1_8001_out0;
wire v_G1_8002_out0;
wire v_G1_8003_out0;
wire v_G1_8004_out0;
wire v_G1_8005_out0;
wire v_G1_8006_out0;
wire v_G1_8007_out0;
wire v_G1_8008_out0;
wire v_G1_8009_out0;
wire v_G1_8010_out0;
wire v_G1_8011_out0;
wire v_G1_8012_out0;
wire v_G1_8013_out0;
wire v_G1_8014_out0;
wire v_G1_8015_out0;
wire v_G1_8016_out0;
wire v_G1_8017_out0;
wire v_G1_8018_out0;
wire v_G1_8019_out0;
wire v_G1_8020_out0;
wire v_G1_8021_out0;
wire v_G1_8022_out0;
wire v_G1_8023_out0;
wire v_G1_8024_out0;
wire v_G1_8025_out0;
wire v_G1_8026_out0;
wire v_G1_8027_out0;
wire v_G1_8028_out0;
wire v_G1_8029_out0;
wire v_G1_8030_out0;
wire v_G1_8031_out0;
wire v_G1_8032_out0;
wire v_G1_8033_out0;
wire v_G1_8034_out0;
wire v_G1_8035_out0;
wire v_G1_8036_out0;
wire v_G1_8037_out0;
wire v_G1_8038_out0;
wire v_G1_8039_out0;
wire v_G1_8040_out0;
wire v_G1_8041_out0;
wire v_G1_8042_out0;
wire v_G1_8043_out0;
wire v_G1_8044_out0;
wire v_G1_8045_out0;
wire v_G1_8046_out0;
wire v_G1_8047_out0;
wire v_G1_8048_out0;
wire v_G1_8049_out0;
wire v_G1_8050_out0;
wire v_G1_8051_out0;
wire v_G1_8052_out0;
wire v_G1_8053_out0;
wire v_G1_8054_out0;
wire v_G1_8055_out0;
wire v_G1_8056_out0;
wire v_G1_8057_out0;
wire v_G1_8058_out0;
wire v_G1_8059_out0;
wire v_G1_8060_out0;
wire v_G1_8061_out0;
wire v_G1_8062_out0;
wire v_G1_8063_out0;
wire v_G1_8064_out0;
wire v_G1_8065_out0;
wire v_G1_8066_out0;
wire v_G1_8067_out0;
wire v_G1_8068_out0;
wire v_G1_8069_out0;
wire v_G1_8070_out0;
wire v_G1_8071_out0;
wire v_G1_8072_out0;
wire v_G1_8073_out0;
wire v_G1_8074_out0;
wire v_G1_8075_out0;
wire v_G1_8076_out0;
wire v_G1_8077_out0;
wire v_G1_8078_out0;
wire v_G1_8079_out0;
wire v_G1_8080_out0;
wire v_G1_8081_out0;
wire v_G1_8082_out0;
wire v_G1_8083_out0;
wire v_G1_8084_out0;
wire v_G1_8085_out0;
wire v_G1_8086_out0;
wire v_G1_8087_out0;
wire v_G1_8088_out0;
wire v_G1_8089_out0;
wire v_G1_8090_out0;
wire v_G1_8091_out0;
wire v_G1_8092_out0;
wire v_G1_8093_out0;
wire v_G1_8094_out0;
wire v_G1_8095_out0;
wire v_G1_8096_out0;
wire v_G1_8097_out0;
wire v_G1_8098_out0;
wire v_G1_8099_out0;
wire v_G1_8100_out0;
wire v_G1_8101_out0;
wire v_G1_8102_out0;
wire v_G1_8103_out0;
wire v_G1_8104_out0;
wire v_G1_8105_out0;
wire v_G1_8106_out0;
wire v_G1_8107_out0;
wire v_G1_8108_out0;
wire v_G1_8109_out0;
wire v_G1_8110_out0;
wire v_G1_8111_out0;
wire v_G1_8112_out0;
wire v_G1_8113_out0;
wire v_G1_8114_out0;
wire v_G1_8115_out0;
wire v_G1_8116_out0;
wire v_G1_8117_out0;
wire v_G1_8118_out0;
wire v_G1_8119_out0;
wire v_G1_8120_out0;
wire v_G1_8121_out0;
wire v_G1_8122_out0;
wire v_G1_8123_out0;
wire v_G1_8124_out0;
wire v_G1_8125_out0;
wire v_G1_8126_out0;
wire v_G1_8127_out0;
wire v_G1_8128_out0;
wire v_G1_8129_out0;
wire v_G1_8130_out0;
wire v_G1_8131_out0;
wire v_G1_8132_out0;
wire v_G1_8133_out0;
wire v_G1_8134_out0;
wire v_G1_8135_out0;
wire v_G1_8136_out0;
wire v_G1_8137_out0;
wire v_G1_8138_out0;
wire v_G1_8139_out0;
wire v_G1_8140_out0;
wire v_G1_8141_out0;
wire v_G1_8142_out0;
wire v_G1_8143_out0;
wire v_G1_8144_out0;
wire v_G1_8145_out0;
wire v_G1_8146_out0;
wire v_G1_8147_out0;
wire v_G1_8148_out0;
wire v_G1_8149_out0;
wire v_G1_8150_out0;
wire v_G1_8151_out0;
wire v_G1_8152_out0;
wire v_G1_8153_out0;
wire v_G1_8154_out0;
wire v_G1_8155_out0;
wire v_G1_8156_out0;
wire v_G1_8157_out0;
wire v_G1_8158_out0;
wire v_G1_8159_out0;
wire v_G1_8160_out0;
wire v_G1_8161_out0;
wire v_G1_8162_out0;
wire v_G1_8163_out0;
wire v_G1_8164_out0;
wire v_G1_8165_out0;
wire v_G1_8166_out0;
wire v_G1_8167_out0;
wire v_G1_8168_out0;
wire v_G1_8169_out0;
wire v_G1_8170_out0;
wire v_G1_8171_out0;
wire v_G1_8172_out0;
wire v_G1_8173_out0;
wire v_G1_8174_out0;
wire v_G1_8175_out0;
wire v_G1_8176_out0;
wire v_G1_8177_out0;
wire v_G1_8178_out0;
wire v_G1_8179_out0;
wire v_G1_8180_out0;
wire v_G1_8181_out0;
wire v_G1_8182_out0;
wire v_G1_8183_out0;
wire v_G1_8184_out0;
wire v_G1_8185_out0;
wire v_G1_8186_out0;
wire v_G1_8187_out0;
wire v_G1_8188_out0;
wire v_G1_8189_out0;
wire v_G1_8190_out0;
wire v_G1_8191_out0;
wire v_G1_8192_out0;
wire v_G1_8193_out0;
wire v_G1_8194_out0;
wire v_G1_8195_out0;
wire v_G1_8196_out0;
wire v_G1_8197_out0;
wire v_G1_8198_out0;
wire v_G1_8199_out0;
wire v_G1_8200_out0;
wire v_G1_8201_out0;
wire v_G1_8202_out0;
wire v_G1_8203_out0;
wire v_G1_8204_out0;
wire v_G1_8205_out0;
wire v_G1_8206_out0;
wire v_G1_8207_out0;
wire v_G1_8208_out0;
wire v_G1_8209_out0;
wire v_G1_8210_out0;
wire v_G1_8211_out0;
wire v_G1_8212_out0;
wire v_G1_8213_out0;
wire v_G1_8214_out0;
wire v_G1_8215_out0;
wire v_G1_8216_out0;
wire v_G1_8217_out0;
wire v_G1_8218_out0;
wire v_G1_8219_out0;
wire v_G1_8220_out0;
wire v_G1_8221_out0;
wire v_G1_8222_out0;
wire v_G1_8223_out0;
wire v_G1_8224_out0;
wire v_G1_8225_out0;
wire v_G1_8226_out0;
wire v_G1_8227_out0;
wire v_G1_8228_out0;
wire v_G1_8229_out0;
wire v_G1_8230_out0;
wire v_G1_8231_out0;
wire v_G1_8232_out0;
wire v_G1_8233_out0;
wire v_G1_8234_out0;
wire v_G1_8235_out0;
wire v_G1_8236_out0;
wire v_G1_8237_out0;
wire v_G1_8238_out0;
wire v_G1_8239_out0;
wire v_G1_8240_out0;
wire v_G1_8241_out0;
wire v_G1_8242_out0;
wire v_G1_8243_out0;
wire v_G1_8244_out0;
wire v_G1_8245_out0;
wire v_G1_8246_out0;
wire v_G1_8247_out0;
wire v_G1_8248_out0;
wire v_G1_8249_out0;
wire v_G1_8250_out0;
wire v_G1_8251_out0;
wire v_G1_8252_out0;
wire v_G1_8253_out0;
wire v_G1_8254_out0;
wire v_G1_8255_out0;
wire v_G1_8256_out0;
wire v_G1_8257_out0;
wire v_G1_8258_out0;
wire v_G1_8259_out0;
wire v_G1_8260_out0;
wire v_G1_8261_out0;
wire v_G1_8262_out0;
wire v_G1_8263_out0;
wire v_G1_8264_out0;
wire v_G1_8265_out0;
wire v_G1_8266_out0;
wire v_G1_8267_out0;
wire v_G1_8268_out0;
wire v_G1_8269_out0;
wire v_G1_8270_out0;
wire v_G1_8271_out0;
wire v_G1_8272_out0;
wire v_G1_8273_out0;
wire v_G1_8274_out0;
wire v_G1_8275_out0;
wire v_G1_8276_out0;
wire v_G1_8277_out0;
wire v_G1_8278_out0;
wire v_G1_8279_out0;
wire v_G1_8280_out0;
wire v_G1_8281_out0;
wire v_G1_8282_out0;
wire v_G1_8283_out0;
wire v_G1_8284_out0;
wire v_G1_8285_out0;
wire v_G1_8286_out0;
wire v_G1_8287_out0;
wire v_G1_8288_out0;
wire v_G1_8289_out0;
wire v_G1_8290_out0;
wire v_G1_8291_out0;
wire v_G1_8292_out0;
wire v_G1_8293_out0;
wire v_G1_8294_out0;
wire v_G1_8295_out0;
wire v_G1_8296_out0;
wire v_G1_8297_out0;
wire v_G1_8298_out0;
wire v_G1_8299_out0;
wire v_G1_8300_out0;
wire v_G1_8301_out0;
wire v_G1_8302_out0;
wire v_G1_8303_out0;
wire v_G1_8304_out0;
wire v_G1_8305_out0;
wire v_G1_8306_out0;
wire v_G1_8307_out0;
wire v_G1_8308_out0;
wire v_G1_8309_out0;
wire v_G1_8310_out0;
wire v_G1_8311_out0;
wire v_G1_8312_out0;
wire v_G1_8313_out0;
wire v_G1_8314_out0;
wire v_G1_8315_out0;
wire v_G1_8316_out0;
wire v_G1_8317_out0;
wire v_G1_8318_out0;
wire v_G1_8319_out0;
wire v_G1_8320_out0;
wire v_G1_8321_out0;
wire v_G1_8322_out0;
wire v_G1_8323_out0;
wire v_G1_8324_out0;
wire v_G1_8325_out0;
wire v_G1_8326_out0;
wire v_G1_8327_out0;
wire v_G1_8328_out0;
wire v_G1_8329_out0;
wire v_G1_8330_out0;
wire v_G1_8331_out0;
wire v_G1_8332_out0;
wire v_G1_8333_out0;
wire v_G1_8334_out0;
wire v_G1_8335_out0;
wire v_G1_8336_out0;
wire v_G1_8337_out0;
wire v_G1_8338_out0;
wire v_G1_8339_out0;
wire v_G1_8340_out0;
wire v_G1_8341_out0;
wire v_G1_8342_out0;
wire v_G1_8343_out0;
wire v_G1_8344_out0;
wire v_G1_8345_out0;
wire v_G1_8346_out0;
wire v_G1_8347_out0;
wire v_G1_8348_out0;
wire v_G1_8349_out0;
wire v_G1_8350_out0;
wire v_G1_8351_out0;
wire v_G1_8352_out0;
wire v_G1_8353_out0;
wire v_G1_8354_out0;
wire v_G1_8355_out0;
wire v_G1_8356_out0;
wire v_G1_8357_out0;
wire v_G1_8358_out0;
wire v_G1_8359_out0;
wire v_G1_8360_out0;
wire v_G1_8361_out0;
wire v_G1_8362_out0;
wire v_G1_8363_out0;
wire v_G1_8364_out0;
wire v_G1_8365_out0;
wire v_G1_8366_out0;
wire v_G1_8367_out0;
wire v_G1_8368_out0;
wire v_G1_8369_out0;
wire v_G1_8370_out0;
wire v_G1_8371_out0;
wire v_G1_8372_out0;
wire v_G1_8373_out0;
wire v_G1_8374_out0;
wire v_G1_8375_out0;
wire v_G1_8376_out0;
wire v_G1_8377_out0;
wire v_G1_8378_out0;
wire v_G1_8379_out0;
wire v_G1_8380_out0;
wire v_G1_8381_out0;
wire v_G1_8382_out0;
wire v_G1_8383_out0;
wire v_G1_8384_out0;
wire v_G1_8385_out0;
wire v_G1_8386_out0;
wire v_G1_8387_out0;
wire v_G1_8388_out0;
wire v_G1_8389_out0;
wire v_G1_8390_out0;
wire v_G1_8391_out0;
wire v_G1_8392_out0;
wire v_G1_8393_out0;
wire v_G1_8394_out0;
wire v_G1_8395_out0;
wire v_G1_8396_out0;
wire v_G1_8397_out0;
wire v_G1_8398_out0;
wire v_G1_8399_out0;
wire v_G1_8400_out0;
wire v_G1_8401_out0;
wire v_G1_8402_out0;
wire v_G1_8403_out0;
wire v_G1_8404_out0;
wire v_G1_8405_out0;
wire v_G1_8406_out0;
wire v_G1_8407_out0;
wire v_G1_8408_out0;
wire v_G1_8409_out0;
wire v_G1_8410_out0;
wire v_G1_8411_out0;
wire v_G1_8412_out0;
wire v_G1_8413_out0;
wire v_G1_8414_out0;
wire v_G1_8415_out0;
wire v_G1_8416_out0;
wire v_G1_8417_out0;
wire v_G1_8418_out0;
wire v_G1_8419_out0;
wire v_G1_8420_out0;
wire v_G1_8421_out0;
wire v_G1_8422_out0;
wire v_G1_8423_out0;
wire v_G1_8424_out0;
wire v_G1_8425_out0;
wire v_G1_8426_out0;
wire v_G1_8427_out0;
wire v_G1_8428_out0;
wire v_G1_8429_out0;
wire v_G1_8430_out0;
wire v_G1_8431_out0;
wire v_G1_8432_out0;
wire v_G1_8433_out0;
wire v_G1_8434_out0;
wire v_G1_8435_out0;
wire v_G1_8436_out0;
wire v_G1_8437_out0;
wire v_G1_8438_out0;
wire v_G1_8439_out0;
wire v_G1_8440_out0;
wire v_G1_8441_out0;
wire v_G1_8442_out0;
wire v_G1_8443_out0;
wire v_G1_8444_out0;
wire v_G1_8445_out0;
wire v_G1_8446_out0;
wire v_G1_8447_out0;
wire v_G1_8448_out0;
wire v_G1_8449_out0;
wire v_G1_8450_out0;
wire v_G1_8451_out0;
wire v_G1_8452_out0;
wire v_G1_8453_out0;
wire v_G1_8454_out0;
wire v_G1_8455_out0;
wire v_G1_8456_out0;
wire v_G1_8457_out0;
wire v_G1_8458_out0;
wire v_G1_8459_out0;
wire v_G1_8460_out0;
wire v_G1_8461_out0;
wire v_G1_8462_out0;
wire v_G1_8463_out0;
wire v_G1_8464_out0;
wire v_G1_8465_out0;
wire v_G1_8466_out0;
wire v_G1_8467_out0;
wire v_G1_8468_out0;
wire v_G1_8469_out0;
wire v_G1_8470_out0;
wire v_G1_8471_out0;
wire v_G1_8472_out0;
wire v_G1_8473_out0;
wire v_G1_8474_out0;
wire v_G1_8475_out0;
wire v_G1_8476_out0;
wire v_G1_8477_out0;
wire v_G1_8478_out0;
wire v_G1_8479_out0;
wire v_G1_8480_out0;
wire v_G1_8481_out0;
wire v_G1_8482_out0;
wire v_G1_8483_out0;
wire v_G1_8484_out0;
wire v_G1_8485_out0;
wire v_G1_8486_out0;
wire v_G1_8487_out0;
wire v_G1_8488_out0;
wire v_G1_8489_out0;
wire v_G1_8490_out0;
wire v_G1_8491_out0;
wire v_G1_8492_out0;
wire v_G1_8493_out0;
wire v_G1_8494_out0;
wire v_G1_8495_out0;
wire v_G1_8496_out0;
wire v_G1_8497_out0;
wire v_G1_8498_out0;
wire v_G1_8499_out0;
wire v_G1_8500_out0;
wire v_G1_8501_out0;
wire v_G1_8502_out0;
wire v_G1_8503_out0;
wire v_G1_8504_out0;
wire v_G1_8505_out0;
wire v_G1_8506_out0;
wire v_G1_8507_out0;
wire v_G1_8508_out0;
wire v_G1_8509_out0;
wire v_G1_8510_out0;
wire v_G1_8511_out0;
wire v_G1_8512_out0;
wire v_G1_8513_out0;
wire v_G1_8514_out0;
wire v_G1_8515_out0;
wire v_G1_8516_out0;
wire v_G1_8517_out0;
wire v_G1_8518_out0;
wire v_G1_8519_out0;
wire v_G1_8520_out0;
wire v_G1_8521_out0;
wire v_G1_8522_out0;
wire v_G1_8523_out0;
wire v_G1_8524_out0;
wire v_G1_8525_out0;
wire v_G1_8526_out0;
wire v_G1_8527_out0;
wire v_G1_8528_out0;
wire v_G1_8529_out0;
wire v_G1_8530_out0;
wire v_G1_8531_out0;
wire v_G1_8532_out0;
wire v_G1_8533_out0;
wire v_G1_8534_out0;
wire v_G1_8535_out0;
wire v_G1_8536_out0;
wire v_G1_8537_out0;
wire v_G1_8538_out0;
wire v_G1_8539_out0;
wire v_G1_8540_out0;
wire v_G1_8541_out0;
wire v_G1_8542_out0;
wire v_G1_8543_out0;
wire v_G1_8544_out0;
wire v_G1_8545_out0;
wire v_G1_8546_out0;
wire v_G1_8547_out0;
wire v_G1_8548_out0;
wire v_G1_8549_out0;
wire v_G1_8550_out0;
wire v_G1_8551_out0;
wire v_G1_8552_out0;
wire v_G1_8553_out0;
wire v_G1_8554_out0;
wire v_G1_8555_out0;
wire v_G1_8556_out0;
wire v_G1_8557_out0;
wire v_G1_8558_out0;
wire v_G1_8559_out0;
wire v_G1_8560_out0;
wire v_G1_8561_out0;
wire v_G1_8562_out0;
wire v_G1_8563_out0;
wire v_G1_8564_out0;
wire v_G1_8565_out0;
wire v_G1_8566_out0;
wire v_G1_8567_out0;
wire v_G1_8568_out0;
wire v_G1_8569_out0;
wire v_G1_8570_out0;
wire v_G1_8571_out0;
wire v_G1_8572_out0;
wire v_G1_8573_out0;
wire v_G1_8574_out0;
wire v_G1_8575_out0;
wire v_G1_8576_out0;
wire v_G1_8577_out0;
wire v_G1_8578_out0;
wire v_G1_8579_out0;
wire v_G1_8580_out0;
wire v_G1_8581_out0;
wire v_G1_8582_out0;
wire v_G1_8583_out0;
wire v_G1_8584_out0;
wire v_G1_8585_out0;
wire v_G1_8586_out0;
wire v_G1_8587_out0;
wire v_G1_8588_out0;
wire v_G1_8589_out0;
wire v_G1_8590_out0;
wire v_G1_8591_out0;
wire v_G1_8592_out0;
wire v_G1_8593_out0;
wire v_G1_8594_out0;
wire v_G1_8595_out0;
wire v_G1_8596_out0;
wire v_G1_8597_out0;
wire v_G1_8598_out0;
wire v_G1_8599_out0;
wire v_G1_8600_out0;
wire v_G1_8601_out0;
wire v_G1_8602_out0;
wire v_G1_8603_out0;
wire v_G1_8604_out0;
wire v_G1_8605_out0;
wire v_G1_8606_out0;
wire v_G1_8607_out0;
wire v_G1_8608_out0;
wire v_G1_8609_out0;
wire v_G1_8610_out0;
wire v_G1_8611_out0;
wire v_G1_8612_out0;
wire v_G1_8613_out0;
wire v_G1_8614_out0;
wire v_G1_8615_out0;
wire v_G1_8616_out0;
wire v_G1_8617_out0;
wire v_G1_8618_out0;
wire v_G1_8619_out0;
wire v_G1_8620_out0;
wire v_G1_8621_out0;
wire v_G1_8622_out0;
wire v_G1_8623_out0;
wire v_G1_8624_out0;
wire v_G1_8625_out0;
wire v_G1_8626_out0;
wire v_G1_8627_out0;
wire v_G1_8628_out0;
wire v_G1_8629_out0;
wire v_G1_8630_out0;
wire v_G1_8631_out0;
wire v_G1_8632_out0;
wire v_G1_8633_out0;
wire v_G1_8634_out0;
wire v_G1_8635_out0;
wire v_G1_8636_out0;
wire v_G1_8637_out0;
wire v_G1_8638_out0;
wire v_G1_8639_out0;
wire v_G1_8640_out0;
wire v_G1_8641_out0;
wire v_G1_8642_out0;
wire v_G1_8643_out0;
wire v_G1_8644_out0;
wire v_G1_8693_out0;
wire v_G1_8694_out0;
wire v_G1_8695_out0;
wire v_G1_8696_out0;
wire v_G20_11040_out0;
wire v_G20_11147_out0;
wire v_G20_11148_out0;
wire v_G20_598_out0;
wire v_G20_599_out0;
wire v_G21_10681_out0;
wire v_G21_10788_out0;
wire v_G21_2656_out0;
wire v_G21_2657_out0;
wire v_G21_2885_out0;
wire v_G21_2886_out0;
wire v_G21_3808_out0;
wire v_G21_3809_out0;
wire v_G21_3810_out0;
wire v_G21_3811_out0;
wire v_G22_10620_out0;
wire v_G22_10983_out0;
wire v_G22_10984_out0;
wire v_G22_10985_out0;
wire v_G22_10986_out0;
wire v_G22_13663_out0;
wire v_G22_13707_out0;
wire v_G22_13708_out0;
wire v_G22_1899_out0;
wire v_G22_1900_out0;
wire v_G23_10439_out0;
wire v_G23_10440_out0;
wire v_G23_2614_out0;
wire v_G23_2840_out0;
wire v_G23_2841_out0;
wire v_G23_3083_out0;
wire v_G23_4852_out0;
wire v_G23_4853_out0;
wire v_G23_4854_out0;
wire v_G23_4855_out0;
wire v_G24_10460_out0;
wire v_G24_10560_out0;
wire v_G24_10561_out0;
wire v_G24_10562_out0;
wire v_G24_10563_out0;
wire v_G24_3955_out0;
wire v_G24_3956_out0;
wire v_G24_4780_out0;
wire v_G25_4658_out0;
wire v_G25_6962_out0;
wire v_G25_6963_out0;
wire v_G26_4735_out0;
wire v_G26_4736_out0;
wire v_G27_9793_out0;
wire v_G27_9794_out0;
wire v_G28_2098_out0;
wire v_G28_2099_out0;
wire v_G28_2100_out0;
wire v_G28_2101_out0;
wire v_G28_6868_out0;
wire v_G28_6869_out0;
wire v_G29_5834_out0;
wire v_G29_5835_out0;
wire v_G2_10278_out0;
wire v_G2_10471_out0;
wire v_G2_10799_out0;
wire v_G2_10800_out0;
wire v_G2_11134_out0;
wire v_G2_11135_out0;
wire v_G2_12230_out0;
wire v_G2_12231_out0;
wire v_G2_12253_out0;
wire v_G2_12254_out0;
wire v_G2_12255_out0;
wire v_G2_12256_out0;
wire v_G2_12257_out0;
wire v_G2_12258_out0;
wire v_G2_12259_out0;
wire v_G2_12260_out0;
wire v_G2_12261_out0;
wire v_G2_12262_out0;
wire v_G2_12263_out0;
wire v_G2_12264_out0;
wire v_G2_12265_out0;
wire v_G2_12266_out0;
wire v_G2_12267_out0;
wire v_G2_12268_out0;
wire v_G2_12269_out0;
wire v_G2_12270_out0;
wire v_G2_12271_out0;
wire v_G2_12272_out0;
wire v_G2_12273_out0;
wire v_G2_12274_out0;
wire v_G2_12275_out0;
wire v_G2_12276_out0;
wire v_G2_12277_out0;
wire v_G2_12278_out0;
wire v_G2_12279_out0;
wire v_G2_12280_out0;
wire v_G2_12281_out0;
wire v_G2_12282_out0;
wire v_G2_12283_out0;
wire v_G2_12284_out0;
wire v_G2_12285_out0;
wire v_G2_12286_out0;
wire v_G2_12287_out0;
wire v_G2_12288_out0;
wire v_G2_12289_out0;
wire v_G2_12290_out0;
wire v_G2_12291_out0;
wire v_G2_12292_out0;
wire v_G2_12293_out0;
wire v_G2_12294_out0;
wire v_G2_12295_out0;
wire v_G2_12296_out0;
wire v_G2_12297_out0;
wire v_G2_12298_out0;
wire v_G2_12299_out0;
wire v_G2_12300_out0;
wire v_G2_12301_out0;
wire v_G2_12302_out0;
wire v_G2_12303_out0;
wire v_G2_12304_out0;
wire v_G2_12305_out0;
wire v_G2_12306_out0;
wire v_G2_12307_out0;
wire v_G2_12308_out0;
wire v_G2_12309_out0;
wire v_G2_12310_out0;
wire v_G2_12311_out0;
wire v_G2_12312_out0;
wire v_G2_12313_out0;
wire v_G2_12314_out0;
wire v_G2_12315_out0;
wire v_G2_12316_out0;
wire v_G2_12317_out0;
wire v_G2_12318_out0;
wire v_G2_12319_out0;
wire v_G2_12320_out0;
wire v_G2_12321_out0;
wire v_G2_12322_out0;
wire v_G2_12323_out0;
wire v_G2_12324_out0;
wire v_G2_12325_out0;
wire v_G2_12326_out0;
wire v_G2_12327_out0;
wire v_G2_12328_out0;
wire v_G2_12329_out0;
wire v_G2_12330_out0;
wire v_G2_12331_out0;
wire v_G2_12332_out0;
wire v_G2_12333_out0;
wire v_G2_12334_out0;
wire v_G2_12335_out0;
wire v_G2_12336_out0;
wire v_G2_12337_out0;
wire v_G2_12338_out0;
wire v_G2_12339_out0;
wire v_G2_12340_out0;
wire v_G2_12341_out0;
wire v_G2_12342_out0;
wire v_G2_12343_out0;
wire v_G2_12344_out0;
wire v_G2_12345_out0;
wire v_G2_12346_out0;
wire v_G2_12347_out0;
wire v_G2_12348_out0;
wire v_G2_12349_out0;
wire v_G2_12350_out0;
wire v_G2_12351_out0;
wire v_G2_12352_out0;
wire v_G2_12353_out0;
wire v_G2_12354_out0;
wire v_G2_12355_out0;
wire v_G2_12356_out0;
wire v_G2_12357_out0;
wire v_G2_12358_out0;
wire v_G2_12359_out0;
wire v_G2_12360_out0;
wire v_G2_12361_out0;
wire v_G2_12362_out0;
wire v_G2_12363_out0;
wire v_G2_12364_out0;
wire v_G2_12365_out0;
wire v_G2_12366_out0;
wire v_G2_12367_out0;
wire v_G2_12368_out0;
wire v_G2_12369_out0;
wire v_G2_12370_out0;
wire v_G2_12371_out0;
wire v_G2_12372_out0;
wire v_G2_12373_out0;
wire v_G2_12374_out0;
wire v_G2_12375_out0;
wire v_G2_12376_out0;
wire v_G2_12377_out0;
wire v_G2_12378_out0;
wire v_G2_12379_out0;
wire v_G2_12380_out0;
wire v_G2_12381_out0;
wire v_G2_12382_out0;
wire v_G2_12383_out0;
wire v_G2_12384_out0;
wire v_G2_12385_out0;
wire v_G2_12386_out0;
wire v_G2_12387_out0;
wire v_G2_12388_out0;
wire v_G2_12389_out0;
wire v_G2_12390_out0;
wire v_G2_12391_out0;
wire v_G2_12392_out0;
wire v_G2_12393_out0;
wire v_G2_12394_out0;
wire v_G2_12395_out0;
wire v_G2_12396_out0;
wire v_G2_12397_out0;
wire v_G2_12398_out0;
wire v_G2_12399_out0;
wire v_G2_12400_out0;
wire v_G2_12401_out0;
wire v_G2_12402_out0;
wire v_G2_12403_out0;
wire v_G2_12404_out0;
wire v_G2_12405_out0;
wire v_G2_12406_out0;
wire v_G2_12407_out0;
wire v_G2_12408_out0;
wire v_G2_12409_out0;
wire v_G2_12410_out0;
wire v_G2_12411_out0;
wire v_G2_12412_out0;
wire v_G2_12413_out0;
wire v_G2_12414_out0;
wire v_G2_12415_out0;
wire v_G2_12416_out0;
wire v_G2_12417_out0;
wire v_G2_12418_out0;
wire v_G2_12419_out0;
wire v_G2_12420_out0;
wire v_G2_12421_out0;
wire v_G2_12422_out0;
wire v_G2_12423_out0;
wire v_G2_12424_out0;
wire v_G2_12425_out0;
wire v_G2_12426_out0;
wire v_G2_12427_out0;
wire v_G2_12428_out0;
wire v_G2_12429_out0;
wire v_G2_12430_out0;
wire v_G2_12431_out0;
wire v_G2_12432_out0;
wire v_G2_12433_out0;
wire v_G2_12434_out0;
wire v_G2_12435_out0;
wire v_G2_12436_out0;
wire v_G2_12437_out0;
wire v_G2_12438_out0;
wire v_G2_12439_out0;
wire v_G2_12440_out0;
wire v_G2_12441_out0;
wire v_G2_12442_out0;
wire v_G2_12443_out0;
wire v_G2_12444_out0;
wire v_G2_12445_out0;
wire v_G2_12446_out0;
wire v_G2_12447_out0;
wire v_G2_12448_out0;
wire v_G2_12449_out0;
wire v_G2_12450_out0;
wire v_G2_12451_out0;
wire v_G2_12452_out0;
wire v_G2_12453_out0;
wire v_G2_12454_out0;
wire v_G2_12455_out0;
wire v_G2_12456_out0;
wire v_G2_12457_out0;
wire v_G2_12458_out0;
wire v_G2_12459_out0;
wire v_G2_12460_out0;
wire v_G2_12461_out0;
wire v_G2_12462_out0;
wire v_G2_12463_out0;
wire v_G2_12464_out0;
wire v_G2_12465_out0;
wire v_G2_12466_out0;
wire v_G2_12467_out0;
wire v_G2_12468_out0;
wire v_G2_12469_out0;
wire v_G2_12470_out0;
wire v_G2_12471_out0;
wire v_G2_12472_out0;
wire v_G2_12473_out0;
wire v_G2_12474_out0;
wire v_G2_12475_out0;
wire v_G2_12476_out0;
wire v_G2_12477_out0;
wire v_G2_12478_out0;
wire v_G2_12479_out0;
wire v_G2_12480_out0;
wire v_G2_12481_out0;
wire v_G2_12482_out0;
wire v_G2_12483_out0;
wire v_G2_12484_out0;
wire v_G2_12485_out0;
wire v_G2_12486_out0;
wire v_G2_12487_out0;
wire v_G2_12488_out0;
wire v_G2_12489_out0;
wire v_G2_12490_out0;
wire v_G2_12491_out0;
wire v_G2_12492_out0;
wire v_G2_12493_out0;
wire v_G2_12494_out0;
wire v_G2_12495_out0;
wire v_G2_12496_out0;
wire v_G2_12497_out0;
wire v_G2_12498_out0;
wire v_G2_12499_out0;
wire v_G2_12500_out0;
wire v_G2_12501_out0;
wire v_G2_12502_out0;
wire v_G2_12503_out0;
wire v_G2_12504_out0;
wire v_G2_12505_out0;
wire v_G2_12506_out0;
wire v_G2_12507_out0;
wire v_G2_12508_out0;
wire v_G2_12509_out0;
wire v_G2_12510_out0;
wire v_G2_12511_out0;
wire v_G2_12512_out0;
wire v_G2_12513_out0;
wire v_G2_12514_out0;
wire v_G2_12515_out0;
wire v_G2_12516_out0;
wire v_G2_12517_out0;
wire v_G2_12518_out0;
wire v_G2_12519_out0;
wire v_G2_12520_out0;
wire v_G2_12521_out0;
wire v_G2_12522_out0;
wire v_G2_12523_out0;
wire v_G2_12524_out0;
wire v_G2_12525_out0;
wire v_G2_12526_out0;
wire v_G2_12527_out0;
wire v_G2_12528_out0;
wire v_G2_12529_out0;
wire v_G2_12530_out0;
wire v_G2_12531_out0;
wire v_G2_12532_out0;
wire v_G2_12533_out0;
wire v_G2_12534_out0;
wire v_G2_12535_out0;
wire v_G2_12536_out0;
wire v_G2_12537_out0;
wire v_G2_12538_out0;
wire v_G2_12539_out0;
wire v_G2_12540_out0;
wire v_G2_12541_out0;
wire v_G2_12542_out0;
wire v_G2_12543_out0;
wire v_G2_12544_out0;
wire v_G2_12545_out0;
wire v_G2_12546_out0;
wire v_G2_12547_out0;
wire v_G2_12548_out0;
wire v_G2_12549_out0;
wire v_G2_12550_out0;
wire v_G2_12551_out0;
wire v_G2_12552_out0;
wire v_G2_12553_out0;
wire v_G2_12554_out0;
wire v_G2_12555_out0;
wire v_G2_12556_out0;
wire v_G2_12557_out0;
wire v_G2_12558_out0;
wire v_G2_12559_out0;
wire v_G2_12560_out0;
wire v_G2_12561_out0;
wire v_G2_12562_out0;
wire v_G2_12563_out0;
wire v_G2_12564_out0;
wire v_G2_12565_out0;
wire v_G2_12566_out0;
wire v_G2_12567_out0;
wire v_G2_12568_out0;
wire v_G2_12569_out0;
wire v_G2_12570_out0;
wire v_G2_12571_out0;
wire v_G2_12572_out0;
wire v_G2_12573_out0;
wire v_G2_12574_out0;
wire v_G2_12575_out0;
wire v_G2_12576_out0;
wire v_G2_12577_out0;
wire v_G2_12578_out0;
wire v_G2_12579_out0;
wire v_G2_12580_out0;
wire v_G2_12581_out0;
wire v_G2_12582_out0;
wire v_G2_12583_out0;
wire v_G2_12584_out0;
wire v_G2_12585_out0;
wire v_G2_12586_out0;
wire v_G2_12587_out0;
wire v_G2_12588_out0;
wire v_G2_12589_out0;
wire v_G2_12590_out0;
wire v_G2_12591_out0;
wire v_G2_12592_out0;
wire v_G2_12593_out0;
wire v_G2_12594_out0;
wire v_G2_12595_out0;
wire v_G2_12596_out0;
wire v_G2_12597_out0;
wire v_G2_12598_out0;
wire v_G2_12599_out0;
wire v_G2_12600_out0;
wire v_G2_12601_out0;
wire v_G2_12602_out0;
wire v_G2_12603_out0;
wire v_G2_12604_out0;
wire v_G2_12605_out0;
wire v_G2_12606_out0;
wire v_G2_12607_out0;
wire v_G2_12608_out0;
wire v_G2_12609_out0;
wire v_G2_12610_out0;
wire v_G2_12611_out0;
wire v_G2_12612_out0;
wire v_G2_12613_out0;
wire v_G2_12614_out0;
wire v_G2_12615_out0;
wire v_G2_12616_out0;
wire v_G2_12617_out0;
wire v_G2_12618_out0;
wire v_G2_12619_out0;
wire v_G2_12620_out0;
wire v_G2_12621_out0;
wire v_G2_12622_out0;
wire v_G2_12623_out0;
wire v_G2_12624_out0;
wire v_G2_12625_out0;
wire v_G2_12626_out0;
wire v_G2_12627_out0;
wire v_G2_12628_out0;
wire v_G2_12629_out0;
wire v_G2_12630_out0;
wire v_G2_12631_out0;
wire v_G2_12632_out0;
wire v_G2_12633_out0;
wire v_G2_12634_out0;
wire v_G2_12635_out0;
wire v_G2_12636_out0;
wire v_G2_12637_out0;
wire v_G2_12638_out0;
wire v_G2_12639_out0;
wire v_G2_12640_out0;
wire v_G2_12641_out0;
wire v_G2_12642_out0;
wire v_G2_12643_out0;
wire v_G2_12644_out0;
wire v_G2_12645_out0;
wire v_G2_12646_out0;
wire v_G2_12647_out0;
wire v_G2_12648_out0;
wire v_G2_12649_out0;
wire v_G2_12650_out0;
wire v_G2_12651_out0;
wire v_G2_12652_out0;
wire v_G2_12653_out0;
wire v_G2_12654_out0;
wire v_G2_12655_out0;
wire v_G2_12656_out0;
wire v_G2_12657_out0;
wire v_G2_12658_out0;
wire v_G2_12659_out0;
wire v_G2_12660_out0;
wire v_G2_12661_out0;
wire v_G2_12662_out0;
wire v_G2_12663_out0;
wire v_G2_12664_out0;
wire v_G2_12665_out0;
wire v_G2_12666_out0;
wire v_G2_12667_out0;
wire v_G2_12668_out0;
wire v_G2_12669_out0;
wire v_G2_12670_out0;
wire v_G2_12671_out0;
wire v_G2_12672_out0;
wire v_G2_12673_out0;
wire v_G2_12674_out0;
wire v_G2_12675_out0;
wire v_G2_12676_out0;
wire v_G2_12677_out0;
wire v_G2_12678_out0;
wire v_G2_12679_out0;
wire v_G2_12680_out0;
wire v_G2_12681_out0;
wire v_G2_12682_out0;
wire v_G2_12683_out0;
wire v_G2_12684_out0;
wire v_G2_12685_out0;
wire v_G2_12686_out0;
wire v_G2_12687_out0;
wire v_G2_12688_out0;
wire v_G2_12689_out0;
wire v_G2_12690_out0;
wire v_G2_12691_out0;
wire v_G2_12692_out0;
wire v_G2_12693_out0;
wire v_G2_12694_out0;
wire v_G2_12695_out0;
wire v_G2_12696_out0;
wire v_G2_12697_out0;
wire v_G2_12698_out0;
wire v_G2_12699_out0;
wire v_G2_12700_out0;
wire v_G2_12701_out0;
wire v_G2_12702_out0;
wire v_G2_12703_out0;
wire v_G2_12704_out0;
wire v_G2_12705_out0;
wire v_G2_12706_out0;
wire v_G2_12707_out0;
wire v_G2_12708_out0;
wire v_G2_12709_out0;
wire v_G2_12710_out0;
wire v_G2_12711_out0;
wire v_G2_12712_out0;
wire v_G2_12713_out0;
wire v_G2_12714_out0;
wire v_G2_12715_out0;
wire v_G2_12716_out0;
wire v_G2_12717_out0;
wire v_G2_12718_out0;
wire v_G2_12719_out0;
wire v_G2_12720_out0;
wire v_G2_12721_out0;
wire v_G2_12722_out0;
wire v_G2_12723_out0;
wire v_G2_12724_out0;
wire v_G2_12725_out0;
wire v_G2_12726_out0;
wire v_G2_12727_out0;
wire v_G2_12728_out0;
wire v_G2_12729_out0;
wire v_G2_12730_out0;
wire v_G2_12731_out0;
wire v_G2_12732_out0;
wire v_G2_12733_out0;
wire v_G2_12734_out0;
wire v_G2_12735_out0;
wire v_G2_12736_out0;
wire v_G2_12737_out0;
wire v_G2_12738_out0;
wire v_G2_12739_out0;
wire v_G2_12740_out0;
wire v_G2_12741_out0;
wire v_G2_12742_out0;
wire v_G2_12743_out0;
wire v_G2_12744_out0;
wire v_G2_12745_out0;
wire v_G2_12746_out0;
wire v_G2_12747_out0;
wire v_G2_12748_out0;
wire v_G2_12749_out0;
wire v_G2_12750_out0;
wire v_G2_12751_out0;
wire v_G2_12752_out0;
wire v_G2_12753_out0;
wire v_G2_12754_out0;
wire v_G2_12755_out0;
wire v_G2_12756_out0;
wire v_G2_12757_out0;
wire v_G2_12758_out0;
wire v_G2_12759_out0;
wire v_G2_12760_out0;
wire v_G2_12761_out0;
wire v_G2_12762_out0;
wire v_G2_12763_out0;
wire v_G2_12764_out0;
wire v_G2_12765_out0;
wire v_G2_12766_out0;
wire v_G2_12767_out0;
wire v_G2_12768_out0;
wire v_G2_12769_out0;
wire v_G2_12770_out0;
wire v_G2_12771_out0;
wire v_G2_12772_out0;
wire v_G2_12773_out0;
wire v_G2_12774_out0;
wire v_G2_12775_out0;
wire v_G2_12776_out0;
wire v_G2_12777_out0;
wire v_G2_12778_out0;
wire v_G2_12779_out0;
wire v_G2_12780_out0;
wire v_G2_12781_out0;
wire v_G2_12782_out0;
wire v_G2_12783_out0;
wire v_G2_12784_out0;
wire v_G2_12785_out0;
wire v_G2_12786_out0;
wire v_G2_12787_out0;
wire v_G2_12788_out0;
wire v_G2_12789_out0;
wire v_G2_12790_out0;
wire v_G2_12791_out0;
wire v_G2_12792_out0;
wire v_G2_12793_out0;
wire v_G2_12794_out0;
wire v_G2_12795_out0;
wire v_G2_12796_out0;
wire v_G2_12797_out0;
wire v_G2_12798_out0;
wire v_G2_12799_out0;
wire v_G2_12800_out0;
wire v_G2_12801_out0;
wire v_G2_12802_out0;
wire v_G2_12803_out0;
wire v_G2_12804_out0;
wire v_G2_12805_out0;
wire v_G2_12806_out0;
wire v_G2_12807_out0;
wire v_G2_12808_out0;
wire v_G2_12809_out0;
wire v_G2_12810_out0;
wire v_G2_12811_out0;
wire v_G2_12812_out0;
wire v_G2_12813_out0;
wire v_G2_12814_out0;
wire v_G2_12815_out0;
wire v_G2_12816_out0;
wire v_G2_12817_out0;
wire v_G2_12818_out0;
wire v_G2_12819_out0;
wire v_G2_12820_out0;
wire v_G2_12821_out0;
wire v_G2_12822_out0;
wire v_G2_12823_out0;
wire v_G2_12824_out0;
wire v_G2_12825_out0;
wire v_G2_12826_out0;
wire v_G2_12827_out0;
wire v_G2_12828_out0;
wire v_G2_12829_out0;
wire v_G2_12830_out0;
wire v_G2_12831_out0;
wire v_G2_12832_out0;
wire v_G2_12833_out0;
wire v_G2_12834_out0;
wire v_G2_12835_out0;
wire v_G2_12836_out0;
wire v_G2_12837_out0;
wire v_G2_12838_out0;
wire v_G2_12839_out0;
wire v_G2_12840_out0;
wire v_G2_12841_out0;
wire v_G2_12842_out0;
wire v_G2_12843_out0;
wire v_G2_12844_out0;
wire v_G2_12845_out0;
wire v_G2_12846_out0;
wire v_G2_12847_out0;
wire v_G2_12848_out0;
wire v_G2_12849_out0;
wire v_G2_12850_out0;
wire v_G2_12851_out0;
wire v_G2_12852_out0;
wire v_G2_12853_out0;
wire v_G2_12854_out0;
wire v_G2_12855_out0;
wire v_G2_12856_out0;
wire v_G2_12857_out0;
wire v_G2_12858_out0;
wire v_G2_12859_out0;
wire v_G2_12860_out0;
wire v_G2_12861_out0;
wire v_G2_12862_out0;
wire v_G2_12863_out0;
wire v_G2_12864_out0;
wire v_G2_12865_out0;
wire v_G2_12866_out0;
wire v_G2_12867_out0;
wire v_G2_12868_out0;
wire v_G2_12869_out0;
wire v_G2_12870_out0;
wire v_G2_12871_out0;
wire v_G2_12872_out0;
wire v_G2_12873_out0;
wire v_G2_12874_out0;
wire v_G2_12875_out0;
wire v_G2_12876_out0;
wire v_G2_12877_out0;
wire v_G2_12878_out0;
wire v_G2_12879_out0;
wire v_G2_12880_out0;
wire v_G2_12881_out0;
wire v_G2_12882_out0;
wire v_G2_12883_out0;
wire v_G2_12884_out0;
wire v_G2_12885_out0;
wire v_G2_12886_out0;
wire v_G2_12887_out0;
wire v_G2_12888_out0;
wire v_G2_12889_out0;
wire v_G2_12890_out0;
wire v_G2_12891_out0;
wire v_G2_12892_out0;
wire v_G2_12893_out0;
wire v_G2_12894_out0;
wire v_G2_12895_out0;
wire v_G2_12896_out0;
wire v_G2_12897_out0;
wire v_G2_12898_out0;
wire v_G2_12899_out0;
wire v_G2_12900_out0;
wire v_G2_12901_out0;
wire v_G2_12902_out0;
wire v_G2_12903_out0;
wire v_G2_12904_out0;
wire v_G2_12905_out0;
wire v_G2_12906_out0;
wire v_G2_12907_out0;
wire v_G2_12908_out0;
wire v_G2_12909_out0;
wire v_G2_12910_out0;
wire v_G2_12911_out0;
wire v_G2_12912_out0;
wire v_G2_12913_out0;
wire v_G2_12914_out0;
wire v_G2_12915_out0;
wire v_G2_12916_out0;
wire v_G2_12917_out0;
wire v_G2_12918_out0;
wire v_G2_12919_out0;
wire v_G2_12920_out0;
wire v_G2_12921_out0;
wire v_G2_12922_out0;
wire v_G2_12923_out0;
wire v_G2_12924_out0;
wire v_G2_12925_out0;
wire v_G2_12926_out0;
wire v_G2_12927_out0;
wire v_G2_12928_out0;
wire v_G2_12929_out0;
wire v_G2_12930_out0;
wire v_G2_12931_out0;
wire v_G2_12932_out0;
wire v_G2_12933_out0;
wire v_G2_12934_out0;
wire v_G2_12935_out0;
wire v_G2_12936_out0;
wire v_G2_12937_out0;
wire v_G2_12938_out0;
wire v_G2_12939_out0;
wire v_G2_12940_out0;
wire v_G2_12941_out0;
wire v_G2_12942_out0;
wire v_G2_12943_out0;
wire v_G2_12944_out0;
wire v_G2_12945_out0;
wire v_G2_12946_out0;
wire v_G2_12947_out0;
wire v_G2_12948_out0;
wire v_G2_12949_out0;
wire v_G2_12950_out0;
wire v_G2_12951_out0;
wire v_G2_12952_out0;
wire v_G2_12953_out0;
wire v_G2_12954_out0;
wire v_G2_12955_out0;
wire v_G2_12956_out0;
wire v_G2_12957_out0;
wire v_G2_12958_out0;
wire v_G2_12959_out0;
wire v_G2_12960_out0;
wire v_G2_12961_out0;
wire v_G2_12962_out0;
wire v_G2_12963_out0;
wire v_G2_12964_out0;
wire v_G2_12965_out0;
wire v_G2_12966_out0;
wire v_G2_12967_out0;
wire v_G2_12968_out0;
wire v_G2_12969_out0;
wire v_G2_12970_out0;
wire v_G2_12971_out0;
wire v_G2_12972_out0;
wire v_G2_12973_out0;
wire v_G2_12974_out0;
wire v_G2_12975_out0;
wire v_G2_12976_out0;
wire v_G2_12977_out0;
wire v_G2_12978_out0;
wire v_G2_12979_out0;
wire v_G2_12980_out0;
wire v_G2_12981_out0;
wire v_G2_12982_out0;
wire v_G2_12983_out0;
wire v_G2_12984_out0;
wire v_G2_12985_out0;
wire v_G2_12986_out0;
wire v_G2_12987_out0;
wire v_G2_12988_out0;
wire v_G2_12989_out0;
wire v_G2_12990_out0;
wire v_G2_12991_out0;
wire v_G2_12992_out0;
wire v_G2_12993_out0;
wire v_G2_12994_out0;
wire v_G2_12995_out0;
wire v_G2_12996_out0;
wire v_G2_12997_out0;
wire v_G2_12998_out0;
wire v_G2_12999_out0;
wire v_G2_13000_out0;
wire v_G2_13001_out0;
wire v_G2_13002_out0;
wire v_G2_13003_out0;
wire v_G2_13004_out0;
wire v_G2_13005_out0;
wire v_G2_13006_out0;
wire v_G2_13007_out0;
wire v_G2_13008_out0;
wire v_G2_13009_out0;
wire v_G2_13010_out0;
wire v_G2_13011_out0;
wire v_G2_13012_out0;
wire v_G2_13013_out0;
wire v_G2_13014_out0;
wire v_G2_13015_out0;
wire v_G2_13016_out0;
wire v_G2_13017_out0;
wire v_G2_13018_out0;
wire v_G2_13019_out0;
wire v_G2_13020_out0;
wire v_G2_13021_out0;
wire v_G2_13022_out0;
wire v_G2_13023_out0;
wire v_G2_13024_out0;
wire v_G2_13025_out0;
wire v_G2_13026_out0;
wire v_G2_13027_out0;
wire v_G2_13028_out0;
wire v_G2_13029_out0;
wire v_G2_13030_out0;
wire v_G2_13031_out0;
wire v_G2_13032_out0;
wire v_G2_13033_out0;
wire v_G2_13034_out0;
wire v_G2_13035_out0;
wire v_G2_13036_out0;
wire v_G2_13037_out0;
wire v_G2_13038_out0;
wire v_G2_13039_out0;
wire v_G2_13040_out0;
wire v_G2_13041_out0;
wire v_G2_13042_out0;
wire v_G2_13043_out0;
wire v_G2_13044_out0;
wire v_G2_13045_out0;
wire v_G2_13046_out0;
wire v_G2_13047_out0;
wire v_G2_13048_out0;
wire v_G2_13049_out0;
wire v_G2_13050_out0;
wire v_G2_13051_out0;
wire v_G2_13052_out0;
wire v_G2_13053_out0;
wire v_G2_13054_out0;
wire v_G2_13055_out0;
wire v_G2_13056_out0;
wire v_G2_13057_out0;
wire v_G2_13058_out0;
wire v_G2_13059_out0;
wire v_G2_13060_out0;
wire v_G2_13061_out0;
wire v_G2_13062_out0;
wire v_G2_13063_out0;
wire v_G2_13064_out0;
wire v_G2_13065_out0;
wire v_G2_13066_out0;
wire v_G2_13067_out0;
wire v_G2_13068_out0;
wire v_G2_13069_out0;
wire v_G2_13070_out0;
wire v_G2_13071_out0;
wire v_G2_13072_out0;
wire v_G2_13073_out0;
wire v_G2_13074_out0;
wire v_G2_13075_out0;
wire v_G2_13076_out0;
wire v_G2_13077_out0;
wire v_G2_13078_out0;
wire v_G2_13079_out0;
wire v_G2_13080_out0;
wire v_G2_13081_out0;
wire v_G2_13082_out0;
wire v_G2_13083_out0;
wire v_G2_13084_out0;
wire v_G2_13085_out0;
wire v_G2_13086_out0;
wire v_G2_13087_out0;
wire v_G2_13088_out0;
wire v_G2_13089_out0;
wire v_G2_13090_out0;
wire v_G2_13091_out0;
wire v_G2_13092_out0;
wire v_G2_13093_out0;
wire v_G2_13094_out0;
wire v_G2_13095_out0;
wire v_G2_13096_out0;
wire v_G2_13097_out0;
wire v_G2_13098_out0;
wire v_G2_13099_out0;
wire v_G2_13100_out0;
wire v_G2_13101_out0;
wire v_G2_13102_out0;
wire v_G2_13103_out0;
wire v_G2_13104_out0;
wire v_G2_13105_out0;
wire v_G2_13106_out0;
wire v_G2_13107_out0;
wire v_G2_13108_out0;
wire v_G2_13109_out0;
wire v_G2_13110_out0;
wire v_G2_13111_out0;
wire v_G2_13112_out0;
wire v_G2_13113_out0;
wire v_G2_13114_out0;
wire v_G2_13115_out0;
wire v_G2_13116_out0;
wire v_G2_13117_out0;
wire v_G2_13118_out0;
wire v_G2_13119_out0;
wire v_G2_13120_out0;
wire v_G2_13121_out0;
wire v_G2_13122_out0;
wire v_G2_13123_out0;
wire v_G2_13124_out0;
wire v_G2_13125_out0;
wire v_G2_13126_out0;
wire v_G2_13127_out0;
wire v_G2_13128_out0;
wire v_G2_13129_out0;
wire v_G2_13130_out0;
wire v_G2_13131_out0;
wire v_G2_13132_out0;
wire v_G2_13133_out0;
wire v_G2_13134_out0;
wire v_G2_13135_out0;
wire v_G2_13136_out0;
wire v_G2_13137_out0;
wire v_G2_13138_out0;
wire v_G2_13139_out0;
wire v_G2_13140_out0;
wire v_G2_13141_out0;
wire v_G2_13142_out0;
wire v_G2_13143_out0;
wire v_G2_13144_out0;
wire v_G2_13145_out0;
wire v_G2_13146_out0;
wire v_G2_13147_out0;
wire v_G2_13148_out0;
wire v_G2_13149_out0;
wire v_G2_13150_out0;
wire v_G2_13151_out0;
wire v_G2_13152_out0;
wire v_G2_13153_out0;
wire v_G2_13154_out0;
wire v_G2_13155_out0;
wire v_G2_13156_out0;
wire v_G2_13157_out0;
wire v_G2_13158_out0;
wire v_G2_13159_out0;
wire v_G2_13160_out0;
wire v_G2_13161_out0;
wire v_G2_13162_out0;
wire v_G2_13163_out0;
wire v_G2_13164_out0;
wire v_G2_13165_out0;
wire v_G2_13166_out0;
wire v_G2_13167_out0;
wire v_G2_13168_out0;
wire v_G2_13169_out0;
wire v_G2_13170_out0;
wire v_G2_13171_out0;
wire v_G2_13172_out0;
wire v_G2_13173_out0;
wire v_G2_13174_out0;
wire v_G2_13175_out0;
wire v_G2_13176_out0;
wire v_G2_13177_out0;
wire v_G2_13178_out0;
wire v_G2_13179_out0;
wire v_G2_13180_out0;
wire v_G2_13645_out0;
wire v_G2_13646_out0;
wire v_G2_1809_out0;
wire v_G2_1810_out0;
wire v_G2_1811_out0;
wire v_G2_1812_out0;
wire v_G2_1887_out0;
wire v_G2_1888_out0;
wire v_G2_2652_out0;
wire v_G2_2653_out0;
wire v_G2_2891_out0;
wire v_G2_2892_out0;
wire v_G2_2975_out0;
wire v_G2_2976_out0;
wire v_G2_2977_out0;
wire v_G2_2978_out0;
wire v_G2_3214_out0;
wire v_G2_3221_out0;
wire v_G2_3239_out0;
wire v_G2_3240_out0;
wire v_G2_3245_out0;
wire v_G2_3246_out0;
wire v_G2_4467_out0;
wire v_G2_4468_out0;
wire v_G2_4620_out0;
wire v_G2_4621_out0;
wire v_G2_4622_out0;
wire v_G2_4623_out0;
wire v_G2_4624_out0;
wire v_G2_4625_out0;
wire v_G2_4626_out0;
wire v_G2_4627_out0;
wire v_G2_4628_out0;
wire v_G2_4629_out0;
wire v_G2_4630_out0;
wire v_G2_4631_out0;
wire v_G2_4632_out0;
wire v_G2_4633_out0;
wire v_G2_4634_out0;
wire v_G2_4635_out0;
wire v_G2_4636_out0;
wire v_G2_4637_out0;
wire v_G2_4638_out0;
wire v_G2_4639_out0;
wire v_G2_4640_out0;
wire v_G2_4641_out0;
wire v_G2_4642_out0;
wire v_G2_4643_out0;
wire v_G2_4644_out0;
wire v_G2_4645_out0;
wire v_G2_4646_out0;
wire v_G2_4647_out0;
wire v_G2_4648_out0;
wire v_G2_4649_out0;
wire v_G2_5840_out0;
wire v_G2_5841_out0;
wire v_G2_6791_out0;
wire v_G2_6792_out0;
wire v_G2_6884_out0;
wire v_G2_6885_out0;
wire v_G2_7015_out0;
wire v_G2_7016_out0;
wire v_G2_7025_out0;
wire v_G2_7026_out0;
wire v_G2_7027_out0;
wire v_G2_7028_out0;
wire v_G30_183_out0;
wire v_G30_184_out0;
wire v_G35_10360_out0;
wire v_G35_10361_out0;
wire v_G35_10362_out0;
wire v_G35_10363_out0;
wire v_G36_3135_out0;
wire v_G36_3136_out0;
wire v_G36_3137_out0;
wire v_G36_3138_out0;
wire v_G37_6900_out0;
wire v_G37_6901_out0;
wire v_G37_6902_out0;
wire v_G37_6903_out0;
wire v_G38_3903_out0;
wire v_G38_3904_out0;
wire v_G38_3905_out0;
wire v_G38_3906_out0;
wire v_G3_10462_out0;
wire v_G3_13507_out0;
wire v_G3_13641_out0;
wire v_G3_13642_out0;
wire v_G3_1720_out0;
wire v_G3_1721_out0;
wire v_G3_17_out0;
wire v_G3_18_out0;
wire v_G3_1949_out0;
wire v_G3_1950_out0;
wire v_G3_206_out0;
wire v_G3_207_out0;
wire v_G3_208_out0;
wire v_G3_209_out0;
wire v_G3_241_out0;
wire v_G3_242_out0;
wire v_G3_243_out0;
wire v_G3_244_out0;
wire v_G3_245_out0;
wire v_G3_246_out0;
wire v_G3_247_out0;
wire v_G3_248_out0;
wire v_G3_249_out0;
wire v_G3_250_out0;
wire v_G3_251_out0;
wire v_G3_252_out0;
wire v_G3_253_out0;
wire v_G3_254_out0;
wire v_G3_255_out0;
wire v_G3_256_out0;
wire v_G3_257_out0;
wire v_G3_258_out0;
wire v_G3_259_out0;
wire v_G3_260_out0;
wire v_G3_261_out0;
wire v_G3_2621_out0;
wire v_G3_2622_out0;
wire v_G3_262_out0;
wire v_G3_263_out0;
wire v_G3_264_out0;
wire v_G3_265_out0;
wire v_G3_266_out0;
wire v_G3_267_out0;
wire v_G3_268_out0;
wire v_G3_2690_out0;
wire v_G3_2691_out0;
wire v_G3_269_out0;
wire v_G3_270_out0;
wire v_G3_2903_out0;
wire v_G3_2904_out0;
wire v_G3_2941_out0;
wire v_G3_2942_out0;
wire v_G3_3343_out0;
wire v_G3_3812_out0;
wire v_G3_3813_out0;
wire v_G3_3948_out0;
wire v_G3_3959_out0;
wire v_G3_3960_out0;
wire v_G3_6894_out0;
wire v_G3_6895_out0;
wire v_G3_6896_out0;
wire v_G3_6897_out0;
wire v_G3_7087_out0;
wire v_G3_7088_out0;
wire v_G3_7089_out0;
wire v_G3_7090_out0;
wire v_G3_8665_out0;
wire v_G3_8666_out0;
wire v_G4_10283_out0;
wire v_G4_10284_out0;
wire v_G4_10997_out0;
wire v_G4_10998_out0;
wire v_G4_10999_out0;
wire v_G4_11000_out0;
wire v_G4_12238_out0;
wire v_G4_12239_out0;
wire v_G4_12243_out0;
wire v_G4_12244_out0;
wire v_G4_13702_out0;
wire v_G4_13703_out0;
wire v_G4_1667_out0;
wire v_G4_1668_out0;
wire v_G4_1960_out0;
wire v_G4_1961_out0;
wire v_G4_1962_out0;
wire v_G4_1963_out0;
wire v_G4_219_out0;
wire v_G4_220_out0;
wire v_G4_2767_out0;
wire v_G4_2768_out0;
wire v_G4_2769_out0;
wire v_G4_2770_out0;
wire v_G4_3235_out0;
wire v_G4_3236_out0;
wire v_G4_341_out0;
wire v_G4_342_out0;
wire v_G4_343_out0;
wire v_G4_344_out0;
wire v_G4_345_out0;
wire v_G4_346_out0;
wire v_G4_347_out0;
wire v_G4_348_out0;
wire v_G4_349_out0;
wire v_G4_350_out0;
wire v_G4_351_out0;
wire v_G4_352_out0;
wire v_G4_353_out0;
wire v_G4_354_out0;
wire v_G4_355_out0;
wire v_G4_356_out0;
wire v_G4_357_out0;
wire v_G4_358_out0;
wire v_G4_359_out0;
wire v_G4_360_out0;
wire v_G4_361_out0;
wire v_G4_362_out0;
wire v_G4_363_out0;
wire v_G4_364_out0;
wire v_G4_365_out0;
wire v_G4_366_out0;
wire v_G4_367_out0;
wire v_G4_368_out0;
wire v_G4_369_out0;
wire v_G4_370_out0;
wire v_G4_381_out0;
wire v_G4_382_out0;
wire v_G4_4738_out0;
wire v_G4_4739_out0;
wire v_G4_4846_out0;
wire v_G4_4847_out0;
wire v_G4_6914_out0;
wire v_G4_6915_out0;
wire v_G5_10441_out0;
wire v_G5_10442_out0;
wire v_G5_10533_out0;
wire v_G5_10534_out0;
wire v_G5_10568_out0;
wire v_G5_10569_out0;
wire v_G5_10570_out0;
wire v_G5_10571_out0;
wire v_G5_10621_out0;
wire v_G5_10622_out0;
wire v_G5_10623_out0;
wire v_G5_10624_out0;
wire v_G5_10625_out0;
wire v_G5_10626_out0;
wire v_G5_10627_out0;
wire v_G5_10628_out0;
wire v_G5_10629_out0;
wire v_G5_10630_out0;
wire v_G5_10631_out0;
wire v_G5_10632_out0;
wire v_G5_10633_out0;
wire v_G5_10634_out0;
wire v_G5_10635_out0;
wire v_G5_10636_out0;
wire v_G5_10637_out0;
wire v_G5_10638_out0;
wire v_G5_10639_out0;
wire v_G5_10640_out0;
wire v_G5_10641_out0;
wire v_G5_10642_out0;
wire v_G5_10643_out0;
wire v_G5_10644_out0;
wire v_G5_10645_out0;
wire v_G5_10646_out0;
wire v_G5_10647_out0;
wire v_G5_10648_out0;
wire v_G5_10649_out0;
wire v_G5_10650_out0;
wire v_G5_10801_out0;
wire v_G5_10914_out0;
wire v_G5_10915_out0;
wire v_G5_10989_out0;
wire v_G5_1198_out0;
wire v_G5_229_out0;
wire v_G5_230_out0;
wire v_G5_2584_out0;
wire v_G5_2585_out0;
wire v_G5_2586_out0;
wire v_G5_2587_out0;
wire v_G5_2756_out0;
wire v_G5_2757_out0;
wire v_G5_2783_out0;
wire v_G5_2784_out0;
wire v_G5_2785_out0;
wire v_G5_2786_out0;
wire v_G5_4477_out0;
wire v_G5_4478_out0;
wire v_G5_454_out0;
wire v_G5_455_out0;
wire v_G5_638_out0;
wire v_G5_639_out0;
wire v_G5_7106_out0;
wire v_G5_7107_out0;
wire v_G6_11143_out0;
wire v_G6_11144_out0;
wire v_G6_1159_out0;
wire v_G6_1160_out0;
wire v_G6_1161_out0;
wire v_G6_1162_out0;
wire v_G6_13258_out0;
wire v_G6_13259_out0;
wire v_G6_13637_out0;
wire v_G6_13638_out0;
wire v_G6_13639_out0;
wire v_G6_13640_out0;
wire v_G6_2116_out0;
wire v_G6_2117_out0;
wire v_G6_2118_out0;
wire v_G6_2119_out0;
wire v_G6_2120_out0;
wire v_G6_2121_out0;
wire v_G6_2122_out0;
wire v_G6_2123_out0;
wire v_G6_2124_out0;
wire v_G6_2125_out0;
wire v_G6_2126_out0;
wire v_G6_2127_out0;
wire v_G6_2128_out0;
wire v_G6_2129_out0;
wire v_G6_2130_out0;
wire v_G6_2131_out0;
wire v_G6_2132_out0;
wire v_G6_2133_out0;
wire v_G6_2134_out0;
wire v_G6_2135_out0;
wire v_G6_2136_out0;
wire v_G6_2137_out0;
wire v_G6_2138_out0;
wire v_G6_2139_out0;
wire v_G6_2140_out0;
wire v_G6_2141_out0;
wire v_G6_2142_out0;
wire v_G6_2143_out0;
wire v_G6_2144_out0;
wire v_G6_2145_out0;
wire v_G6_2416_out0;
wire v_G6_2417_out0;
wire v_G6_2905_out0;
wire v_G6_2906_out0;
wire v_G6_327_out0;
wire v_G6_328_out0;
wire v_G6_4531_out0;
wire v_G6_4818_out0;
wire v_G6_8834_out0;
wire v_G6_8835_out0;
wire v_G6_8836_out0;
wire v_G6_8837_out0;
wire v_G7_10332_out0;
wire v_G7_11095_out0;
wire v_G7_11262_out0;
wire v_G7_11263_out0;
wire v_G7_11264_out0;
wire v_G7_11265_out0;
wire v_G7_11266_out0;
wire v_G7_11267_out0;
wire v_G7_11268_out0;
wire v_G7_11269_out0;
wire v_G7_11270_out0;
wire v_G7_11271_out0;
wire v_G7_11272_out0;
wire v_G7_11273_out0;
wire v_G7_11274_out0;
wire v_G7_11275_out0;
wire v_G7_11276_out0;
wire v_G7_11277_out0;
wire v_G7_11278_out0;
wire v_G7_11279_out0;
wire v_G7_11280_out0;
wire v_G7_11281_out0;
wire v_G7_11282_out0;
wire v_G7_11283_out0;
wire v_G7_11284_out0;
wire v_G7_11285_out0;
wire v_G7_11286_out0;
wire v_G7_11287_out0;
wire v_G7_11288_out0;
wire v_G7_11289_out0;
wire v_G7_11290_out0;
wire v_G7_11291_out0;
wire v_G7_1197_out0;
wire v_G7_1684_out0;
wire v_G7_1685_out0;
wire v_G7_169_out0;
wire v_G7_170_out0;
wire v_G7_2455_out0;
wire v_G7_2779_out0;
wire v_G7_2780_out0;
wire v_G7_2781_out0;
wire v_G7_2782_out0;
wire v_G7_4474_out0;
wire v_G7_4475_out0;
wire v_G7_4821_out0;
wire v_G7_4822_out0;
wire v_G7_6862_out0;
wire v_G7_6863_out0;
wire v_G7_8655_out0;
wire v_G7_8656_out0;
wire v_G7_8657_out0;
wire v_G7_8658_out0;
wire v_G8_10609_out0;
wire v_G8_10610_out0;
wire v_G8_10611_out0;
wire v_G8_10612_out0;
wire v_G8_10769_out0;
wire v_G8_10770_out0;
wire v_G8_1215_out0;
wire v_G8_1216_out0;
wire v_G8_1217_out0;
wire v_G8_1218_out0;
wire v_G8_16_out0;
wire v_G8_1765_out0;
wire v_G8_1766_out0;
wire v_G8_2024_out0;
wire v_G8_2025_out0;
wire v_G8_2472_out0;
wire v_G8_2473_out0;
wire v_G8_2474_out0;
wire v_G8_2475_out0;
wire v_G8_2476_out0;
wire v_G8_2477_out0;
wire v_G8_2478_out0;
wire v_G8_2479_out0;
wire v_G8_2480_out0;
wire v_G8_2481_out0;
wire v_G8_2482_out0;
wire v_G8_2483_out0;
wire v_G8_2484_out0;
wire v_G8_2485_out0;
wire v_G8_2486_out0;
wire v_G8_2487_out0;
wire v_G8_2488_out0;
wire v_G8_2489_out0;
wire v_G8_2490_out0;
wire v_G8_2491_out0;
wire v_G8_2492_out0;
wire v_G8_2493_out0;
wire v_G8_2494_out0;
wire v_G8_2495_out0;
wire v_G8_2496_out0;
wire v_G8_2497_out0;
wire v_G8_2498_out0;
wire v_G8_2499_out0;
wire v_G8_2500_out0;
wire v_G8_2501_out0;
wire v_G8_2623_out0;
wire v_G8_2624_out0;
wire v_G8_2644_out0;
wire v_G8_4453_out0;
wire v_G8_4454_out0;
wire v_G8_548_out0;
wire v_G8_549_out0;
wire v_G8_550_out0;
wire v_G8_551_out0;
wire v_G8_7103_out0;
wire v_G9_10291_out0;
wire v_G9_10292_out0;
wire v_G9_10293_out0;
wire v_G9_10294_out0;
wire v_G9_10572_out0;
wire v_G9_10573_out0;
wire v_G9_10574_out0;
wire v_G9_10575_out0;
wire v_G9_10576_out0;
wire v_G9_10577_out0;
wire v_G9_10578_out0;
wire v_G9_10579_out0;
wire v_G9_10580_out0;
wire v_G9_10581_out0;
wire v_G9_10582_out0;
wire v_G9_10583_out0;
wire v_G9_10584_out0;
wire v_G9_10585_out0;
wire v_G9_10586_out0;
wire v_G9_10587_out0;
wire v_G9_10588_out0;
wire v_G9_10589_out0;
wire v_G9_10590_out0;
wire v_G9_10591_out0;
wire v_G9_10592_out0;
wire v_G9_10593_out0;
wire v_G9_10594_out0;
wire v_G9_10595_out0;
wire v_G9_10596_out0;
wire v_G9_10597_out0;
wire v_G9_10598_out0;
wire v_G9_10599_out0;
wire v_G9_10600_out0;
wire v_G9_10601_out0;
wire v_G9_13285_out0;
wire v_G9_13286_out0;
wire v_G9_13287_out0;
wire v_G9_13288_out0;
wire v_G9_13340_out0;
wire v_G9_13341_out0;
wire v_G9_13564_out0;
wire v_G9_13655_out0;
wire v_G9_1671_out0;
wire v_G9_1672_out0;
wire v_G9_223_out0;
wire v_G9_2332_out0;
wire v_G9_2333_out0;
wire v_G9_2895_out0;
wire v_G9_2896_out0;
wire v_G9_2897_out0;
wire v_G9_2898_out0;
wire v_G9_407_out0;
wire v_G9_408_out0;
wire v_G9_411_out0;
wire v_G9_412_out0;
wire v_IN_2466_out0;
wire v_IR15_2464_out0;
wire v_IR15_2465_out0;
wire v_JEQZ_10514_out0;
wire v_JEQZ_10515_out0;
wire v_JEQZ_2981_out0;
wire v_JEQZ_2982_out0;
wire v_JEQ_10496_out0;
wire v_JEQ_10497_out0;
wire v_JEQ_13560_out0;
wire v_JEQ_13561_out0;
wire v_JEQ_2234_out0;
wire v_JEQ_2235_out0;
wire v_JEQ_4445_out0;
wire v_JEQ_4446_out0;
wire v_JEQ_8806_out0;
wire v_JEQ_8807_out0;
wire v_JMIN_1205_out0;
wire v_JMIN_1206_out0;
wire v_JMIN_2662_out0;
wire v_JMIN_2663_out0;
wire v_JMI_13349_out0;
wire v_JMI_13350_out0;
wire v_JMI_1939_out0;
wire v_JMI_1940_out0;
wire v_JMI_3212_out0;
wire v_JMI_3213_out0;
wire v_JMI_8679_out0;
wire v_JMI_8680_out0;
wire v_JMI_88_out0;
wire v_JMI_89_out0;
wire v_JMP_2668_out0;
wire v_JMP_2669_out0;
wire v_JMP_3233_out0;
wire v_JMP_3234_out0;
wire v_JMP_546_out0;
wire v_JMP_547_out0;
wire v_JMP_7077_out0;
wire v_JMP_7078_out0;
wire v_JMP_8825_out0;
wire v_JMP_8826_out0;
wire v_JUMP_2187_out0;
wire v_JUMP_2188_out0;
wire v_LDR_STR0_10349_out0;
wire v_LDR_STR1_13616_out0;
wire v_LOAD_231_out0;
wire v_LOAD_232_out0;
wire v_LOAD_2899_out0;
wire v_LOAD_2900_out0;
wire v_LOAD_3115_out0;
wire v_LOAD_3116_out0;
wire v_LOAD_3949_out0;
wire v_LOAD_3950_out0;
wire v_LOAD_7110_out0;
wire v_LOAD_7111_out0;
wire v_LOAD_8765_out0;
wire v_LOAD_8766_out0;
wire v_LS0_4548_out0;
wire v_LS1_3169_out0;
wire v_LSL_1861_out0;
wire v_LSL_1862_out0;
wire v_LSL_2842_out0;
wire v_LSL_2843_out0;
wire v_LSL_3047_out0;
wire v_LSL_3048_out0;
wire v_LSL_3182_out0;
wire v_LSL_3183_out0;
wire v_LSR_1174_out0;
wire v_LSR_1175_out0;
wire v_LSR_13331_out0;
wire v_LSR_13332_out0;
wire v_LSR_418_out0;
wire v_LSR_419_out0;
wire v_LSR_6912_out0;
wire v_LSR_6913_out0;
wire v_LS_1202_out0;
wire v_LS_1203_out0;
wire v_LS_202_out0;
wire v_LS_203_out0;
wire v_LS_204_out0;
wire v_LS_205_out0;
wire v_LS_2864_out0;
wire v_LS_2865_out0;
wire v_MI_10833_out0;
wire v_MI_10834_out0;
wire v_MI_2612_out0;
wire v_MI_2613_out0;
wire v_MI_560_out0;
wire v_MI_561_out0;
wire v_MOV_10389_out0;
wire v_MOV_10390_out0;
wire v_MOV_196_out0;
wire v_MOV_197_out0;
wire v_MULTI_INSTRUCTION_13308_out0;
wire v_MULTI_INSTRUCTION_13309_out0;
wire v_MULTI_INSTRUCTION_13323_out0;
wire v_MULTI_INSTRUCTION_13324_out0;
wire v_MULTI_INSTRUCTION_2451_out0;
wire v_MULTI_INSTRUCTION_2452_out0;
wire v_MULTI_INSTRUCTION_3953_out0;
wire v_MULTI_INSTRUCTION_3954_out0;
wire v_MULTI_INSTRUCTION_619_out0;
wire v_MULTI_INSTRUCTION_620_out0;
wire v_MULTI_OPCODE_10797_out0;
wire v_MULTI_OPCODE_10798_out0;
wire v_MULTI_OPCODE_11096_out0;
wire v_MULTI_OPCODE_11097_out0;
wire v_MULTI_OPCODE_3020_out0;
wire v_MULTI_OPCODE_3021_out0;
wire v_MUX1_2625_out0;
wire v_MUX1_650_out0;
wire v_MUX2_1180_out0;
wire v_MUX2_4448_out0;
wire v_MUX3_10994_out0;
wire v_MUX3_7140_out0;
wire v_MUX3_8817_out0;
wire v_MUX3_8818_out0;
wire v_MUX4_3219_out0;
wire v_MUX5_10260_out0;
wire v_MUX5_10261_out0;
wire v_MUX5_13348_out0;
wire v_MUX5_7678_out0;
wire v_MUX6_10976_out0;
wire v_MUX6_8757_out0;
wire v_MUX6_8758_out0;
wire v_MUX7_10448_out0;
wire v_MUX8_2697_out0;
wire v_MUX9_166_out0;
wire v_MUX_ENABLE_2349_out0;
wire v_NEGATIVE_11256_out0;
wire v_NEGATIVE_11257_out0;
wire v_NORMAL0_2307_out0;
wire v_NORMAL1_6790_out0;
wire v_NORMAL_10256_out0;
wire v_NORMAL_10257_out0;
wire v_NORMAL_13429_out0;
wire v_NORMAL_13430_out0;
wire v_NORMAL_181_out0;
wire v_NORMAL_182_out0;
wire v_NORMAL_3353_out0;
wire v_NORMAL_3354_out0;
wire v_NORMAL_7114_out0;
wire v_NORMAL_7115_out0;
wire v_NOTUSED1_10684_out0;
wire v_NOTUSED1_10685_out0;
wire v_NOTUSED2_5794_out0;
wire v_NOTUSED2_5795_out0;
wire v_NOTUSED3_10550_out0;
wire v_NOTUSED3_10551_out0;
wire v_NOTUSED4_10530_out0;
wire v_NOTUSED4_10531_out0;
wire v_NOTUSED_10835_out0;
wire v_NOTUSED_10836_out0;
wire v_NOTUSED_1968_out0;
wire v_NOTUSED_1969_out0;
wire v_NOTUSED_325_out0;
wire v_NOTUSED_326_out0;
wire v_NOTUSED_4463_out0;
wire v_NOTUSED_4464_out0;
wire v_NOTUSED_4609_out0;
wire v_OP2_SIGN_10839_out0;
wire v_OP2_SIGN_10840_out0;
wire v_OP2_SIGN_11208_out0;
wire v_OP2_SIGN_11209_out0;
wire v_OUTSTREAM_2097_out0;
wire v_OUT_22_out0;
wire v_OVERFLOW_10492_out0;
wire v_OVERFLOW_10493_out0;
wire v_P_10682_out0;
wire v_P_10683_out0;
wire v_Q0_11198_out0;
wire v_Q0_11199_out0;
wire v_Q0_11200_out0;
wire v_Q0_11201_out0;
wire v_Q0_13351_out0;
wire v_Q0_4470_out0;
wire v_Q0_4471_out0;
wire v_Q0_4472_out0;
wire v_Q0_4473_out0;
wire v_Q0_625_out0;
wire v_Q0_626_out0;
wire v_Q1_2112_out0;
wire v_Q1_307_out0;
wire v_Q1_308_out0;
wire v_Q1_3993_out0;
wire v_Q1_6906_out0;
wire v_Q1_6907_out0;
wire v_Q1_6908_out0;
wire v_Q1_6909_out0;
wire v_Q1_8859_out0;
wire v_Q1_8860_out0;
wire v_Q1_8861_out0;
wire v_Q1_8862_out0;
wire v_Q2_1676_out0;
wire v_Q2_1677_out0;
wire v_Q2_1678_out0;
wire v_Q2_1679_out0;
wire v_Q2_6880_out0;
wire v_Q2_6881_out0;
wire v_Q2_6882_out0;
wire v_Q2_6883_out0;
wire v_Q3_10518_out0;
wire v_Q3_10519_out0;
wire v_Q3_10520_out0;
wire v_Q3_10521_out0;
wire v_Q3_8737_out0;
wire v_Q3_8738_out0;
wire v_Q3_8739_out0;
wire v_Q3_8740_out0;
wire v_Q6_1889_out0;
wire v_Q6_1890_out0;
wire v_Q6_1891_out0;
wire v_Q6_1892_out0;
wire v_Q7_6888_out0;
wire v_Q7_6889_out0;
wire v_Q7_6890_out0;
wire v_Q7_6891_out0;
wire v_Q_291_out0;
wire v_Q_292_out0;
wire v_Q_293_out0;
wire v_Q_294_out0;
wire v_Q_295_out0;
wire v_Q_296_out0;
wire v_Q_297_out0;
wire v_Q_298_out0;
wire v_Q_299_out0;
wire v_Q_300_out0;
wire v_Q_301_out0;
wire v_Q_302_out0;
wire v_Q_303_out0;
wire v_Q_304_out0;
wire v_Q_305_out0;
wire v_Q_306_out0;
wire v_RAMWEN_10701_out0;
wire v_RAMWEN_10702_out0;
wire v_RDN_3349_out0;
wire v_RDN_3351_out0;
wire v_RDN_4496_out0;
wire v_RDN_4497_out0;
wire v_RDN_4498_out0;
wire v_RDN_4499_out0;
wire v_RDN_4500_out0;
wire v_RDN_4501_out0;
wire v_RDN_4502_out0;
wire v_RDN_4503_out0;
wire v_RDN_4504_out0;
wire v_RDN_4505_out0;
wire v_RDN_4506_out0;
wire v_RDN_4507_out0;
wire v_RDN_4508_out0;
wire v_RDN_4509_out0;
wire v_RDN_4510_out0;
wire v_RDN_4511_out0;
wire v_RDN_4512_out0;
wire v_RDN_4513_out0;
wire v_RDN_4514_out0;
wire v_RDN_4515_out0;
wire v_RDN_4516_out0;
wire v_RDN_4517_out0;
wire v_RDN_4518_out0;
wire v_RDN_4519_out0;
wire v_RDN_4520_out0;
wire v_RDN_4521_out0;
wire v_RDN_4522_out0;
wire v_RDN_4523_out0;
wire v_RDN_4524_out0;
wire v_RDN_4525_out0;
wire v_RD_13567_out0;
wire v_RD_13568_out0;
wire v_RD_13569_out0;
wire v_RD_13570_out0;
wire v_RD_13571_out0;
wire v_RD_13572_out0;
wire v_RD_13573_out0;
wire v_RD_13574_out0;
wire v_RD_13575_out0;
wire v_RD_13576_out0;
wire v_RD_13577_out0;
wire v_RD_13578_out0;
wire v_RD_13579_out0;
wire v_RD_13580_out0;
wire v_RD_13581_out0;
wire v_RD_13582_out0;
wire v_RD_13583_out0;
wire v_RD_13584_out0;
wire v_RD_13585_out0;
wire v_RD_13586_out0;
wire v_RD_13587_out0;
wire v_RD_13588_out0;
wire v_RD_13589_out0;
wire v_RD_13590_out0;
wire v_RD_13591_out0;
wire v_RD_13592_out0;
wire v_RD_13593_out0;
wire v_RD_13594_out0;
wire v_RD_13595_out0;
wire v_RD_13596_out0;
wire v_RD_5862_out0;
wire v_RD_5863_out0;
wire v_RD_5864_out0;
wire v_RD_5865_out0;
wire v_RD_5866_out0;
wire v_RD_5867_out0;
wire v_RD_5868_out0;
wire v_RD_5869_out0;
wire v_RD_5870_out0;
wire v_RD_5871_out0;
wire v_RD_5872_out0;
wire v_RD_5873_out0;
wire v_RD_5874_out0;
wire v_RD_5875_out0;
wire v_RD_5876_out0;
wire v_RD_5877_out0;
wire v_RD_5878_out0;
wire v_RD_5879_out0;
wire v_RD_5880_out0;
wire v_RD_5881_out0;
wire v_RD_5882_out0;
wire v_RD_5883_out0;
wire v_RD_5884_out0;
wire v_RD_5885_out0;
wire v_RD_5886_out0;
wire v_RD_5887_out0;
wire v_RD_5888_out0;
wire v_RD_5889_out0;
wire v_RD_5890_out0;
wire v_RD_5891_out0;
wire v_RD_5892_out0;
wire v_RD_5893_out0;
wire v_RD_5894_out0;
wire v_RD_5895_out0;
wire v_RD_5896_out0;
wire v_RD_5897_out0;
wire v_RD_5898_out0;
wire v_RD_5899_out0;
wire v_RD_5900_out0;
wire v_RD_5901_out0;
wire v_RD_5902_out0;
wire v_RD_5903_out0;
wire v_RD_5904_out0;
wire v_RD_5905_out0;
wire v_RD_5906_out0;
wire v_RD_5907_out0;
wire v_RD_5908_out0;
wire v_RD_5909_out0;
wire v_RD_5910_out0;
wire v_RD_5911_out0;
wire v_RD_5912_out0;
wire v_RD_5913_out0;
wire v_RD_5914_out0;
wire v_RD_5915_out0;
wire v_RD_5916_out0;
wire v_RD_5917_out0;
wire v_RD_5918_out0;
wire v_RD_5919_out0;
wire v_RD_5920_out0;
wire v_RD_5921_out0;
wire v_RD_5922_out0;
wire v_RD_5923_out0;
wire v_RD_5924_out0;
wire v_RD_5925_out0;
wire v_RD_5926_out0;
wire v_RD_5927_out0;
wire v_RD_5928_out0;
wire v_RD_5929_out0;
wire v_RD_5930_out0;
wire v_RD_5931_out0;
wire v_RD_5932_out0;
wire v_RD_5933_out0;
wire v_RD_5934_out0;
wire v_RD_5935_out0;
wire v_RD_5936_out0;
wire v_RD_5937_out0;
wire v_RD_5938_out0;
wire v_RD_5939_out0;
wire v_RD_5940_out0;
wire v_RD_5941_out0;
wire v_RD_5942_out0;
wire v_RD_5943_out0;
wire v_RD_5944_out0;
wire v_RD_5945_out0;
wire v_RD_5946_out0;
wire v_RD_5947_out0;
wire v_RD_5948_out0;
wire v_RD_5949_out0;
wire v_RD_5950_out0;
wire v_RD_5951_out0;
wire v_RD_5952_out0;
wire v_RD_5953_out0;
wire v_RD_5954_out0;
wire v_RD_5955_out0;
wire v_RD_5956_out0;
wire v_RD_5957_out0;
wire v_RD_5958_out0;
wire v_RD_5959_out0;
wire v_RD_5960_out0;
wire v_RD_5961_out0;
wire v_RD_5962_out0;
wire v_RD_5963_out0;
wire v_RD_5964_out0;
wire v_RD_5965_out0;
wire v_RD_5966_out0;
wire v_RD_5967_out0;
wire v_RD_5968_out0;
wire v_RD_5969_out0;
wire v_RD_5970_out0;
wire v_RD_5971_out0;
wire v_RD_5972_out0;
wire v_RD_5973_out0;
wire v_RD_5974_out0;
wire v_RD_5975_out0;
wire v_RD_5976_out0;
wire v_RD_5977_out0;
wire v_RD_5978_out0;
wire v_RD_5979_out0;
wire v_RD_5980_out0;
wire v_RD_5981_out0;
wire v_RD_5982_out0;
wire v_RD_5983_out0;
wire v_RD_5984_out0;
wire v_RD_5985_out0;
wire v_RD_5986_out0;
wire v_RD_5987_out0;
wire v_RD_5988_out0;
wire v_RD_5989_out0;
wire v_RD_5990_out0;
wire v_RD_5991_out0;
wire v_RD_5992_out0;
wire v_RD_5993_out0;
wire v_RD_5994_out0;
wire v_RD_5995_out0;
wire v_RD_5996_out0;
wire v_RD_5997_out0;
wire v_RD_5998_out0;
wire v_RD_5999_out0;
wire v_RD_6000_out0;
wire v_RD_6001_out0;
wire v_RD_6002_out0;
wire v_RD_6003_out0;
wire v_RD_6004_out0;
wire v_RD_6005_out0;
wire v_RD_6006_out0;
wire v_RD_6007_out0;
wire v_RD_6008_out0;
wire v_RD_6009_out0;
wire v_RD_6010_out0;
wire v_RD_6011_out0;
wire v_RD_6012_out0;
wire v_RD_6013_out0;
wire v_RD_6014_out0;
wire v_RD_6015_out0;
wire v_RD_6016_out0;
wire v_RD_6017_out0;
wire v_RD_6018_out0;
wire v_RD_6019_out0;
wire v_RD_6020_out0;
wire v_RD_6021_out0;
wire v_RD_6022_out0;
wire v_RD_6023_out0;
wire v_RD_6024_out0;
wire v_RD_6025_out0;
wire v_RD_6026_out0;
wire v_RD_6027_out0;
wire v_RD_6028_out0;
wire v_RD_6029_out0;
wire v_RD_6030_out0;
wire v_RD_6031_out0;
wire v_RD_6032_out0;
wire v_RD_6033_out0;
wire v_RD_6034_out0;
wire v_RD_6035_out0;
wire v_RD_6036_out0;
wire v_RD_6037_out0;
wire v_RD_6038_out0;
wire v_RD_6039_out0;
wire v_RD_6040_out0;
wire v_RD_6041_out0;
wire v_RD_6042_out0;
wire v_RD_6043_out0;
wire v_RD_6044_out0;
wire v_RD_6045_out0;
wire v_RD_6046_out0;
wire v_RD_6047_out0;
wire v_RD_6048_out0;
wire v_RD_6049_out0;
wire v_RD_6050_out0;
wire v_RD_6051_out0;
wire v_RD_6052_out0;
wire v_RD_6053_out0;
wire v_RD_6054_out0;
wire v_RD_6055_out0;
wire v_RD_6056_out0;
wire v_RD_6057_out0;
wire v_RD_6058_out0;
wire v_RD_6059_out0;
wire v_RD_6060_out0;
wire v_RD_6061_out0;
wire v_RD_6062_out0;
wire v_RD_6063_out0;
wire v_RD_6064_out0;
wire v_RD_6065_out0;
wire v_RD_6066_out0;
wire v_RD_6067_out0;
wire v_RD_6068_out0;
wire v_RD_6069_out0;
wire v_RD_6070_out0;
wire v_RD_6071_out0;
wire v_RD_6072_out0;
wire v_RD_6073_out0;
wire v_RD_6074_out0;
wire v_RD_6075_out0;
wire v_RD_6076_out0;
wire v_RD_6077_out0;
wire v_RD_6078_out0;
wire v_RD_6079_out0;
wire v_RD_6080_out0;
wire v_RD_6081_out0;
wire v_RD_6082_out0;
wire v_RD_6083_out0;
wire v_RD_6084_out0;
wire v_RD_6085_out0;
wire v_RD_6086_out0;
wire v_RD_6087_out0;
wire v_RD_6088_out0;
wire v_RD_6089_out0;
wire v_RD_6090_out0;
wire v_RD_6091_out0;
wire v_RD_6092_out0;
wire v_RD_6093_out0;
wire v_RD_6094_out0;
wire v_RD_6095_out0;
wire v_RD_6096_out0;
wire v_RD_6097_out0;
wire v_RD_6098_out0;
wire v_RD_6099_out0;
wire v_RD_6100_out0;
wire v_RD_6101_out0;
wire v_RD_6102_out0;
wire v_RD_6103_out0;
wire v_RD_6104_out0;
wire v_RD_6105_out0;
wire v_RD_6106_out0;
wire v_RD_6107_out0;
wire v_RD_6108_out0;
wire v_RD_6109_out0;
wire v_RD_6110_out0;
wire v_RD_6111_out0;
wire v_RD_6112_out0;
wire v_RD_6113_out0;
wire v_RD_6114_out0;
wire v_RD_6115_out0;
wire v_RD_6116_out0;
wire v_RD_6117_out0;
wire v_RD_6118_out0;
wire v_RD_6119_out0;
wire v_RD_6120_out0;
wire v_RD_6121_out0;
wire v_RD_6122_out0;
wire v_RD_6123_out0;
wire v_RD_6124_out0;
wire v_RD_6125_out0;
wire v_RD_6126_out0;
wire v_RD_6127_out0;
wire v_RD_6128_out0;
wire v_RD_6129_out0;
wire v_RD_6130_out0;
wire v_RD_6131_out0;
wire v_RD_6132_out0;
wire v_RD_6133_out0;
wire v_RD_6134_out0;
wire v_RD_6135_out0;
wire v_RD_6136_out0;
wire v_RD_6137_out0;
wire v_RD_6138_out0;
wire v_RD_6139_out0;
wire v_RD_6140_out0;
wire v_RD_6141_out0;
wire v_RD_6142_out0;
wire v_RD_6143_out0;
wire v_RD_6144_out0;
wire v_RD_6145_out0;
wire v_RD_6146_out0;
wire v_RD_6147_out0;
wire v_RD_6148_out0;
wire v_RD_6149_out0;
wire v_RD_6150_out0;
wire v_RD_6151_out0;
wire v_RD_6152_out0;
wire v_RD_6153_out0;
wire v_RD_6154_out0;
wire v_RD_6155_out0;
wire v_RD_6156_out0;
wire v_RD_6157_out0;
wire v_RD_6158_out0;
wire v_RD_6159_out0;
wire v_RD_6160_out0;
wire v_RD_6161_out0;
wire v_RD_6162_out0;
wire v_RD_6163_out0;
wire v_RD_6164_out0;
wire v_RD_6165_out0;
wire v_RD_6166_out0;
wire v_RD_6167_out0;
wire v_RD_6168_out0;
wire v_RD_6169_out0;
wire v_RD_6170_out0;
wire v_RD_6171_out0;
wire v_RD_6172_out0;
wire v_RD_6173_out0;
wire v_RD_6174_out0;
wire v_RD_6175_out0;
wire v_RD_6176_out0;
wire v_RD_6177_out0;
wire v_RD_6178_out0;
wire v_RD_6179_out0;
wire v_RD_6180_out0;
wire v_RD_6181_out0;
wire v_RD_6182_out0;
wire v_RD_6183_out0;
wire v_RD_6184_out0;
wire v_RD_6185_out0;
wire v_RD_6186_out0;
wire v_RD_6187_out0;
wire v_RD_6188_out0;
wire v_RD_6189_out0;
wire v_RD_6190_out0;
wire v_RD_6191_out0;
wire v_RD_6192_out0;
wire v_RD_6193_out0;
wire v_RD_6194_out0;
wire v_RD_6195_out0;
wire v_RD_6196_out0;
wire v_RD_6197_out0;
wire v_RD_6198_out0;
wire v_RD_6199_out0;
wire v_RD_6200_out0;
wire v_RD_6201_out0;
wire v_RD_6202_out0;
wire v_RD_6203_out0;
wire v_RD_6204_out0;
wire v_RD_6205_out0;
wire v_RD_6206_out0;
wire v_RD_6207_out0;
wire v_RD_6208_out0;
wire v_RD_6209_out0;
wire v_RD_6210_out0;
wire v_RD_6211_out0;
wire v_RD_6212_out0;
wire v_RD_6213_out0;
wire v_RD_6214_out0;
wire v_RD_6215_out0;
wire v_RD_6216_out0;
wire v_RD_6217_out0;
wire v_RD_6218_out0;
wire v_RD_6219_out0;
wire v_RD_6220_out0;
wire v_RD_6221_out0;
wire v_RD_6222_out0;
wire v_RD_6223_out0;
wire v_RD_6224_out0;
wire v_RD_6225_out0;
wire v_RD_6226_out0;
wire v_RD_6227_out0;
wire v_RD_6228_out0;
wire v_RD_6229_out0;
wire v_RD_6230_out0;
wire v_RD_6231_out0;
wire v_RD_6232_out0;
wire v_RD_6233_out0;
wire v_RD_6234_out0;
wire v_RD_6235_out0;
wire v_RD_6236_out0;
wire v_RD_6237_out0;
wire v_RD_6238_out0;
wire v_RD_6239_out0;
wire v_RD_6240_out0;
wire v_RD_6241_out0;
wire v_RD_6242_out0;
wire v_RD_6243_out0;
wire v_RD_6244_out0;
wire v_RD_6245_out0;
wire v_RD_6246_out0;
wire v_RD_6247_out0;
wire v_RD_6248_out0;
wire v_RD_6249_out0;
wire v_RD_6250_out0;
wire v_RD_6251_out0;
wire v_RD_6252_out0;
wire v_RD_6253_out0;
wire v_RD_6254_out0;
wire v_RD_6255_out0;
wire v_RD_6256_out0;
wire v_RD_6257_out0;
wire v_RD_6258_out0;
wire v_RD_6259_out0;
wire v_RD_6260_out0;
wire v_RD_6261_out0;
wire v_RD_6262_out0;
wire v_RD_6263_out0;
wire v_RD_6264_out0;
wire v_RD_6265_out0;
wire v_RD_6266_out0;
wire v_RD_6267_out0;
wire v_RD_6268_out0;
wire v_RD_6269_out0;
wire v_RD_6270_out0;
wire v_RD_6271_out0;
wire v_RD_6272_out0;
wire v_RD_6273_out0;
wire v_RD_6274_out0;
wire v_RD_6275_out0;
wire v_RD_6276_out0;
wire v_RD_6277_out0;
wire v_RD_6278_out0;
wire v_RD_6279_out0;
wire v_RD_6280_out0;
wire v_RD_6281_out0;
wire v_RD_6282_out0;
wire v_RD_6283_out0;
wire v_RD_6284_out0;
wire v_RD_6285_out0;
wire v_RD_6286_out0;
wire v_RD_6287_out0;
wire v_RD_6288_out0;
wire v_RD_6289_out0;
wire v_RD_6290_out0;
wire v_RD_6291_out0;
wire v_RD_6292_out0;
wire v_RD_6293_out0;
wire v_RD_6294_out0;
wire v_RD_6295_out0;
wire v_RD_6296_out0;
wire v_RD_6297_out0;
wire v_RD_6298_out0;
wire v_RD_6299_out0;
wire v_RD_6300_out0;
wire v_RD_6301_out0;
wire v_RD_6302_out0;
wire v_RD_6303_out0;
wire v_RD_6304_out0;
wire v_RD_6305_out0;
wire v_RD_6306_out0;
wire v_RD_6307_out0;
wire v_RD_6308_out0;
wire v_RD_6309_out0;
wire v_RD_6310_out0;
wire v_RD_6311_out0;
wire v_RD_6312_out0;
wire v_RD_6313_out0;
wire v_RD_6314_out0;
wire v_RD_6315_out0;
wire v_RD_6316_out0;
wire v_RD_6317_out0;
wire v_RD_6318_out0;
wire v_RD_6319_out0;
wire v_RD_6320_out0;
wire v_RD_6321_out0;
wire v_RD_6322_out0;
wire v_RD_6323_out0;
wire v_RD_6324_out0;
wire v_RD_6325_out0;
wire v_RD_6326_out0;
wire v_RD_6327_out0;
wire v_RD_6328_out0;
wire v_RD_6329_out0;
wire v_RD_6330_out0;
wire v_RD_6331_out0;
wire v_RD_6332_out0;
wire v_RD_6333_out0;
wire v_RD_6334_out0;
wire v_RD_6335_out0;
wire v_RD_6336_out0;
wire v_RD_6337_out0;
wire v_RD_6338_out0;
wire v_RD_6339_out0;
wire v_RD_6340_out0;
wire v_RD_6341_out0;
wire v_RD_6342_out0;
wire v_RD_6343_out0;
wire v_RD_6344_out0;
wire v_RD_6345_out0;
wire v_RD_6346_out0;
wire v_RD_6347_out0;
wire v_RD_6348_out0;
wire v_RD_6349_out0;
wire v_RD_6350_out0;
wire v_RD_6351_out0;
wire v_RD_6352_out0;
wire v_RD_6353_out0;
wire v_RD_6354_out0;
wire v_RD_6355_out0;
wire v_RD_6356_out0;
wire v_RD_6357_out0;
wire v_RD_6358_out0;
wire v_RD_6359_out0;
wire v_RD_6360_out0;
wire v_RD_6361_out0;
wire v_RD_6362_out0;
wire v_RD_6363_out0;
wire v_RD_6364_out0;
wire v_RD_6365_out0;
wire v_RD_6366_out0;
wire v_RD_6367_out0;
wire v_RD_6368_out0;
wire v_RD_6369_out0;
wire v_RD_6370_out0;
wire v_RD_6371_out0;
wire v_RD_6372_out0;
wire v_RD_6373_out0;
wire v_RD_6374_out0;
wire v_RD_6375_out0;
wire v_RD_6376_out0;
wire v_RD_6377_out0;
wire v_RD_6378_out0;
wire v_RD_6379_out0;
wire v_RD_6380_out0;
wire v_RD_6381_out0;
wire v_RD_6382_out0;
wire v_RD_6383_out0;
wire v_RD_6384_out0;
wire v_RD_6385_out0;
wire v_RD_6386_out0;
wire v_RD_6387_out0;
wire v_RD_6388_out0;
wire v_RD_6389_out0;
wire v_RD_6390_out0;
wire v_RD_6391_out0;
wire v_RD_6392_out0;
wire v_RD_6393_out0;
wire v_RD_6394_out0;
wire v_RD_6395_out0;
wire v_RD_6396_out0;
wire v_RD_6397_out0;
wire v_RD_6398_out0;
wire v_RD_6399_out0;
wire v_RD_6400_out0;
wire v_RD_6401_out0;
wire v_RD_6402_out0;
wire v_RD_6403_out0;
wire v_RD_6404_out0;
wire v_RD_6405_out0;
wire v_RD_6406_out0;
wire v_RD_6407_out0;
wire v_RD_6408_out0;
wire v_RD_6409_out0;
wire v_RD_6410_out0;
wire v_RD_6411_out0;
wire v_RD_6412_out0;
wire v_RD_6413_out0;
wire v_RD_6414_out0;
wire v_RD_6415_out0;
wire v_RD_6416_out0;
wire v_RD_6417_out0;
wire v_RD_6418_out0;
wire v_RD_6419_out0;
wire v_RD_6420_out0;
wire v_RD_6421_out0;
wire v_RD_6422_out0;
wire v_RD_6423_out0;
wire v_RD_6424_out0;
wire v_RD_6425_out0;
wire v_RD_6426_out0;
wire v_RD_6427_out0;
wire v_RD_6428_out0;
wire v_RD_6429_out0;
wire v_RD_6430_out0;
wire v_RD_6431_out0;
wire v_RD_6432_out0;
wire v_RD_6433_out0;
wire v_RD_6434_out0;
wire v_RD_6435_out0;
wire v_RD_6436_out0;
wire v_RD_6437_out0;
wire v_RD_6438_out0;
wire v_RD_6439_out0;
wire v_RD_6440_out0;
wire v_RD_6441_out0;
wire v_RD_6442_out0;
wire v_RD_6443_out0;
wire v_RD_6444_out0;
wire v_RD_6445_out0;
wire v_RD_6446_out0;
wire v_RD_6447_out0;
wire v_RD_6448_out0;
wire v_RD_6449_out0;
wire v_RD_6450_out0;
wire v_RD_6451_out0;
wire v_RD_6452_out0;
wire v_RD_6453_out0;
wire v_RD_6454_out0;
wire v_RD_6455_out0;
wire v_RD_6456_out0;
wire v_RD_6457_out0;
wire v_RD_6458_out0;
wire v_RD_6459_out0;
wire v_RD_6460_out0;
wire v_RD_6461_out0;
wire v_RD_6462_out0;
wire v_RD_6463_out0;
wire v_RD_6464_out0;
wire v_RD_6465_out0;
wire v_RD_6466_out0;
wire v_RD_6467_out0;
wire v_RD_6468_out0;
wire v_RD_6469_out0;
wire v_RD_6470_out0;
wire v_RD_6471_out0;
wire v_RD_6472_out0;
wire v_RD_6473_out0;
wire v_RD_6474_out0;
wire v_RD_6475_out0;
wire v_RD_6476_out0;
wire v_RD_6477_out0;
wire v_RD_6478_out0;
wire v_RD_6479_out0;
wire v_RD_6480_out0;
wire v_RD_6481_out0;
wire v_RD_6482_out0;
wire v_RD_6483_out0;
wire v_RD_6484_out0;
wire v_RD_6485_out0;
wire v_RD_6486_out0;
wire v_RD_6487_out0;
wire v_RD_6488_out0;
wire v_RD_6489_out0;
wire v_RD_6490_out0;
wire v_RD_6491_out0;
wire v_RD_6492_out0;
wire v_RD_6493_out0;
wire v_RD_6494_out0;
wire v_RD_6495_out0;
wire v_RD_6496_out0;
wire v_RD_6497_out0;
wire v_RD_6498_out0;
wire v_RD_6499_out0;
wire v_RD_6500_out0;
wire v_RD_6501_out0;
wire v_RD_6502_out0;
wire v_RD_6503_out0;
wire v_RD_6504_out0;
wire v_RD_6505_out0;
wire v_RD_6506_out0;
wire v_RD_6507_out0;
wire v_RD_6508_out0;
wire v_RD_6509_out0;
wire v_RD_6510_out0;
wire v_RD_6511_out0;
wire v_RD_6512_out0;
wire v_RD_6513_out0;
wire v_RD_6514_out0;
wire v_RD_6515_out0;
wire v_RD_6516_out0;
wire v_RD_6517_out0;
wire v_RD_6518_out0;
wire v_RD_6519_out0;
wire v_RD_6520_out0;
wire v_RD_6521_out0;
wire v_RD_6522_out0;
wire v_RD_6523_out0;
wire v_RD_6524_out0;
wire v_RD_6525_out0;
wire v_RD_6526_out0;
wire v_RD_6527_out0;
wire v_RD_6528_out0;
wire v_RD_6529_out0;
wire v_RD_6530_out0;
wire v_RD_6531_out0;
wire v_RD_6532_out0;
wire v_RD_6533_out0;
wire v_RD_6534_out0;
wire v_RD_6535_out0;
wire v_RD_6536_out0;
wire v_RD_6537_out0;
wire v_RD_6538_out0;
wire v_RD_6539_out0;
wire v_RD_6540_out0;
wire v_RD_6541_out0;
wire v_RD_6542_out0;
wire v_RD_6543_out0;
wire v_RD_6544_out0;
wire v_RD_6545_out0;
wire v_RD_6546_out0;
wire v_RD_6547_out0;
wire v_RD_6548_out0;
wire v_RD_6549_out0;
wire v_RD_6550_out0;
wire v_RD_6551_out0;
wire v_RD_6552_out0;
wire v_RD_6553_out0;
wire v_RD_6554_out0;
wire v_RD_6555_out0;
wire v_RD_6556_out0;
wire v_RD_6557_out0;
wire v_RD_6558_out0;
wire v_RD_6559_out0;
wire v_RD_6560_out0;
wire v_RD_6561_out0;
wire v_RD_6562_out0;
wire v_RD_6563_out0;
wire v_RD_6564_out0;
wire v_RD_6565_out0;
wire v_RD_6566_out0;
wire v_RD_6567_out0;
wire v_RD_6568_out0;
wire v_RD_6569_out0;
wire v_RD_6570_out0;
wire v_RD_6571_out0;
wire v_RD_6572_out0;
wire v_RD_6573_out0;
wire v_RD_6574_out0;
wire v_RD_6575_out0;
wire v_RD_6576_out0;
wire v_RD_6577_out0;
wire v_RD_6578_out0;
wire v_RD_6579_out0;
wire v_RD_6580_out0;
wire v_RD_6581_out0;
wire v_RD_6582_out0;
wire v_RD_6583_out0;
wire v_RD_6584_out0;
wire v_RD_6585_out0;
wire v_RD_6586_out0;
wire v_RD_6587_out0;
wire v_RD_6588_out0;
wire v_RD_6589_out0;
wire v_RD_6590_out0;
wire v_RD_6591_out0;
wire v_RD_6592_out0;
wire v_RD_6593_out0;
wire v_RD_6594_out0;
wire v_RD_6595_out0;
wire v_RD_6596_out0;
wire v_RD_6597_out0;
wire v_RD_6598_out0;
wire v_RD_6599_out0;
wire v_RD_6600_out0;
wire v_RD_6601_out0;
wire v_RD_6602_out0;
wire v_RD_6603_out0;
wire v_RD_6604_out0;
wire v_RD_6605_out0;
wire v_RD_6606_out0;
wire v_RD_6607_out0;
wire v_RD_6608_out0;
wire v_RD_6609_out0;
wire v_RD_6610_out0;
wire v_RD_6611_out0;
wire v_RD_6612_out0;
wire v_RD_6613_out0;
wire v_RD_6614_out0;
wire v_RD_6615_out0;
wire v_RD_6616_out0;
wire v_RD_6617_out0;
wire v_RD_6618_out0;
wire v_RD_6619_out0;
wire v_RD_6620_out0;
wire v_RD_6621_out0;
wire v_RD_6622_out0;
wire v_RD_6623_out0;
wire v_RD_6624_out0;
wire v_RD_6625_out0;
wire v_RD_6626_out0;
wire v_RD_6627_out0;
wire v_RD_6628_out0;
wire v_RD_6629_out0;
wire v_RD_6630_out0;
wire v_RD_6631_out0;
wire v_RD_6632_out0;
wire v_RD_6633_out0;
wire v_RD_6634_out0;
wire v_RD_6635_out0;
wire v_RD_6636_out0;
wire v_RD_6637_out0;
wire v_RD_6638_out0;
wire v_RD_6639_out0;
wire v_RD_6640_out0;
wire v_RD_6641_out0;
wire v_RD_6642_out0;
wire v_RD_6643_out0;
wire v_RD_6644_out0;
wire v_RD_6645_out0;
wire v_RD_6646_out0;
wire v_RD_6647_out0;
wire v_RD_6648_out0;
wire v_RD_6649_out0;
wire v_RD_6650_out0;
wire v_RD_6651_out0;
wire v_RD_6652_out0;
wire v_RD_6653_out0;
wire v_RD_6654_out0;
wire v_RD_6655_out0;
wire v_RD_6656_out0;
wire v_RD_6657_out0;
wire v_RD_6658_out0;
wire v_RD_6659_out0;
wire v_RD_6660_out0;
wire v_RD_6661_out0;
wire v_RD_6662_out0;
wire v_RD_6663_out0;
wire v_RD_6664_out0;
wire v_RD_6665_out0;
wire v_RD_6666_out0;
wire v_RD_6667_out0;
wire v_RD_6668_out0;
wire v_RD_6669_out0;
wire v_RD_6670_out0;
wire v_RD_6671_out0;
wire v_RD_6672_out0;
wire v_RD_6673_out0;
wire v_RD_6674_out0;
wire v_RD_6675_out0;
wire v_RD_6676_out0;
wire v_RD_6677_out0;
wire v_RD_6678_out0;
wire v_RD_6679_out0;
wire v_RD_6680_out0;
wire v_RD_6681_out0;
wire v_RD_6682_out0;
wire v_RD_6683_out0;
wire v_RD_6684_out0;
wire v_RD_6685_out0;
wire v_RD_6686_out0;
wire v_RD_6687_out0;
wire v_RD_6688_out0;
wire v_RD_6689_out0;
wire v_RD_6690_out0;
wire v_RD_6691_out0;
wire v_RD_6692_out0;
wire v_RD_6693_out0;
wire v_RD_6694_out0;
wire v_RD_6695_out0;
wire v_RD_6696_out0;
wire v_RD_6697_out0;
wire v_RD_6698_out0;
wire v_RD_6699_out0;
wire v_RD_6700_out0;
wire v_RD_6701_out0;
wire v_RD_6702_out0;
wire v_RD_6703_out0;
wire v_RD_6704_out0;
wire v_RD_6705_out0;
wire v_RD_6706_out0;
wire v_RD_6707_out0;
wire v_RD_6708_out0;
wire v_RD_6709_out0;
wire v_RD_6710_out0;
wire v_RD_6711_out0;
wire v_RD_6712_out0;
wire v_RD_6713_out0;
wire v_RD_6714_out0;
wire v_RD_6715_out0;
wire v_RD_6716_out0;
wire v_RD_6717_out0;
wire v_RD_6718_out0;
wire v_RD_6719_out0;
wire v_RD_6720_out0;
wire v_RD_6721_out0;
wire v_RD_6722_out0;
wire v_RD_6723_out0;
wire v_RD_6724_out0;
wire v_RD_6725_out0;
wire v_RD_6726_out0;
wire v_RD_6727_out0;
wire v_RD_6728_out0;
wire v_RD_6729_out0;
wire v_RD_6730_out0;
wire v_RD_6731_out0;
wire v_RD_6732_out0;
wire v_RD_6733_out0;
wire v_RD_6734_out0;
wire v_RD_6735_out0;
wire v_RD_6736_out0;
wire v_RD_6737_out0;
wire v_RD_6738_out0;
wire v_RD_6739_out0;
wire v_RD_6740_out0;
wire v_RD_6741_out0;
wire v_RD_6742_out0;
wire v_RD_6743_out0;
wire v_RD_6744_out0;
wire v_RD_6745_out0;
wire v_RD_6746_out0;
wire v_RD_6747_out0;
wire v_RD_6748_out0;
wire v_RD_6749_out0;
wire v_RD_6750_out0;
wire v_RD_6751_out0;
wire v_RD_6752_out0;
wire v_RD_6753_out0;
wire v_RD_6754_out0;
wire v_RD_6755_out0;
wire v_RD_6756_out0;
wire v_RD_6757_out0;
wire v_RD_6758_out0;
wire v_RD_6759_out0;
wire v_RD_6760_out0;
wire v_RD_6761_out0;
wire v_RD_6762_out0;
wire v_RD_6763_out0;
wire v_RD_6764_out0;
wire v_RD_6765_out0;
wire v_RD_6766_out0;
wire v_RD_6767_out0;
wire v_RD_6768_out0;
wire v_RD_6769_out0;
wire v_RD_6770_out0;
wire v_RD_6771_out0;
wire v_RD_6772_out0;
wire v_RD_6773_out0;
wire v_RD_6774_out0;
wire v_RD_6775_out0;
wire v_RD_6776_out0;
wire v_RD_6777_out0;
wire v_RD_6778_out0;
wire v_RD_6779_out0;
wire v_RD_6780_out0;
wire v_RD_6781_out0;
wire v_RD_6782_out0;
wire v_RD_6783_out0;
wire v_RD_6784_out0;
wire v_RD_6785_out0;
wire v_RD_6786_out0;
wire v_RD_6787_out0;
wire v_RD_6788_out0;
wire v_RD_6789_out0;
wire v_RD_7187_out0;
wire v_RD_7188_out0;
wire v_RD_7189_out0;
wire v_RD_7190_out0;
wire v_RD_7191_out0;
wire v_RD_7192_out0;
wire v_RD_7193_out0;
wire v_RD_7194_out0;
wire v_RD_7195_out0;
wire v_RD_7196_out0;
wire v_RD_7197_out0;
wire v_RD_7198_out0;
wire v_RD_7199_out0;
wire v_RD_7200_out0;
wire v_RD_7201_out0;
wire v_RD_7202_out0;
wire v_RD_7203_out0;
wire v_RD_7204_out0;
wire v_RD_7205_out0;
wire v_RD_7206_out0;
wire v_RD_7207_out0;
wire v_RD_7208_out0;
wire v_RD_7209_out0;
wire v_RD_7210_out0;
wire v_RD_7211_out0;
wire v_RD_7212_out0;
wire v_RD_7213_out0;
wire v_RD_7214_out0;
wire v_RD_7215_out0;
wire v_RD_7216_out0;
wire v_RD_7217_out0;
wire v_RD_7218_out0;
wire v_RD_7219_out0;
wire v_RD_7220_out0;
wire v_RD_7221_out0;
wire v_RD_7222_out0;
wire v_RD_7223_out0;
wire v_RD_7224_out0;
wire v_RD_7225_out0;
wire v_RD_7226_out0;
wire v_RD_7227_out0;
wire v_RD_7228_out0;
wire v_RD_7229_out0;
wire v_RD_7230_out0;
wire v_RD_7231_out0;
wire v_RD_7232_out0;
wire v_RD_7233_out0;
wire v_RD_7234_out0;
wire v_RD_7235_out0;
wire v_RD_7236_out0;
wire v_RD_7237_out0;
wire v_RD_7238_out0;
wire v_RD_7239_out0;
wire v_RD_7240_out0;
wire v_RD_7241_out0;
wire v_RD_7242_out0;
wire v_RD_7243_out0;
wire v_RD_7244_out0;
wire v_RD_7245_out0;
wire v_RD_7246_out0;
wire v_RD_7247_out0;
wire v_RD_7248_out0;
wire v_RD_7249_out0;
wire v_RD_7250_out0;
wire v_RD_7251_out0;
wire v_RD_7252_out0;
wire v_RD_7253_out0;
wire v_RD_7254_out0;
wire v_RD_7255_out0;
wire v_RD_7256_out0;
wire v_RD_7257_out0;
wire v_RD_7258_out0;
wire v_RD_7259_out0;
wire v_RD_7260_out0;
wire v_RD_7261_out0;
wire v_RD_7262_out0;
wire v_RD_7263_out0;
wire v_RD_7264_out0;
wire v_RD_7265_out0;
wire v_RD_7266_out0;
wire v_RD_7267_out0;
wire v_RD_7268_out0;
wire v_RD_7269_out0;
wire v_RD_7270_out0;
wire v_RD_7271_out0;
wire v_RD_7272_out0;
wire v_RD_7273_out0;
wire v_RD_7274_out0;
wire v_RD_7275_out0;
wire v_RD_7276_out0;
wire v_RD_7277_out0;
wire v_RD_7278_out0;
wire v_RD_7279_out0;
wire v_RD_7280_out0;
wire v_RD_7281_out0;
wire v_RD_7282_out0;
wire v_RD_7283_out0;
wire v_RD_7284_out0;
wire v_RD_7285_out0;
wire v_RD_7286_out0;
wire v_RD_7287_out0;
wire v_RD_7288_out0;
wire v_RD_7289_out0;
wire v_RD_7290_out0;
wire v_RD_7291_out0;
wire v_RD_7292_out0;
wire v_RD_7293_out0;
wire v_RD_7294_out0;
wire v_RD_7295_out0;
wire v_RD_7296_out0;
wire v_RD_7297_out0;
wire v_RD_7298_out0;
wire v_RD_7299_out0;
wire v_RD_7300_out0;
wire v_RD_7301_out0;
wire v_RD_7302_out0;
wire v_RD_7303_out0;
wire v_RD_7304_out0;
wire v_RD_7305_out0;
wire v_RD_7306_out0;
wire v_RD_7307_out0;
wire v_RD_7308_out0;
wire v_RD_7309_out0;
wire v_RD_7310_out0;
wire v_RD_7311_out0;
wire v_RD_7312_out0;
wire v_RD_7313_out0;
wire v_RD_7314_out0;
wire v_RD_7315_out0;
wire v_RD_7316_out0;
wire v_RD_7317_out0;
wire v_RD_7318_out0;
wire v_RD_7319_out0;
wire v_RD_7320_out0;
wire v_RD_7321_out0;
wire v_RD_7322_out0;
wire v_RD_7323_out0;
wire v_RD_7324_out0;
wire v_RD_7325_out0;
wire v_RD_7326_out0;
wire v_RD_7327_out0;
wire v_RD_7328_out0;
wire v_RD_7329_out0;
wire v_RD_7330_out0;
wire v_RD_7331_out0;
wire v_RD_7332_out0;
wire v_RD_7333_out0;
wire v_RD_7334_out0;
wire v_RD_7335_out0;
wire v_RD_7336_out0;
wire v_RD_7337_out0;
wire v_RD_7338_out0;
wire v_RD_7339_out0;
wire v_RD_7340_out0;
wire v_RD_7341_out0;
wire v_RD_7342_out0;
wire v_RD_7343_out0;
wire v_RD_7344_out0;
wire v_RD_7345_out0;
wire v_RD_7346_out0;
wire v_RD_7347_out0;
wire v_RD_7348_out0;
wire v_RD_7349_out0;
wire v_RD_7350_out0;
wire v_RD_7351_out0;
wire v_RD_7352_out0;
wire v_RD_7353_out0;
wire v_RD_7354_out0;
wire v_RD_7355_out0;
wire v_RD_7356_out0;
wire v_RD_7357_out0;
wire v_RD_7358_out0;
wire v_RD_7359_out0;
wire v_RD_7360_out0;
wire v_RD_7361_out0;
wire v_RD_7362_out0;
wire v_RD_7363_out0;
wire v_RD_7364_out0;
wire v_RD_7365_out0;
wire v_RD_7366_out0;
wire v_RD_7367_out0;
wire v_RD_7368_out0;
wire v_RD_7369_out0;
wire v_RD_7370_out0;
wire v_RD_7371_out0;
wire v_RD_7372_out0;
wire v_RD_7373_out0;
wire v_RD_7374_out0;
wire v_RD_7375_out0;
wire v_RD_7376_out0;
wire v_RD_7377_out0;
wire v_RD_7378_out0;
wire v_RD_7379_out0;
wire v_RD_7380_out0;
wire v_RD_7381_out0;
wire v_RD_7382_out0;
wire v_RD_7383_out0;
wire v_RD_7384_out0;
wire v_RD_7385_out0;
wire v_RD_7386_out0;
wire v_RD_7387_out0;
wire v_RD_7388_out0;
wire v_RD_7389_out0;
wire v_RD_7390_out0;
wire v_RD_7391_out0;
wire v_RD_7392_out0;
wire v_RD_7393_out0;
wire v_RD_7394_out0;
wire v_RD_7395_out0;
wire v_RD_7396_out0;
wire v_RD_7397_out0;
wire v_RD_7398_out0;
wire v_RD_7399_out0;
wire v_RD_7400_out0;
wire v_RD_7401_out0;
wire v_RD_7402_out0;
wire v_RD_7403_out0;
wire v_RD_7404_out0;
wire v_RD_7405_out0;
wire v_RD_7406_out0;
wire v_RD_7407_out0;
wire v_RD_7408_out0;
wire v_RD_7409_out0;
wire v_RD_7410_out0;
wire v_RD_7411_out0;
wire v_RD_7412_out0;
wire v_RD_7413_out0;
wire v_RD_7414_out0;
wire v_RD_7415_out0;
wire v_RD_7416_out0;
wire v_RD_7417_out0;
wire v_RD_7418_out0;
wire v_RD_7419_out0;
wire v_RD_7420_out0;
wire v_RD_7421_out0;
wire v_RD_7422_out0;
wire v_RD_7423_out0;
wire v_RD_7424_out0;
wire v_RD_7425_out0;
wire v_RD_7426_out0;
wire v_RD_7427_out0;
wire v_RD_7428_out0;
wire v_RD_7429_out0;
wire v_RD_7430_out0;
wire v_RD_7431_out0;
wire v_RD_7432_out0;
wire v_RD_7433_out0;
wire v_RD_7434_out0;
wire v_RD_7435_out0;
wire v_RD_7436_out0;
wire v_RD_7437_out0;
wire v_RD_7438_out0;
wire v_RD_7439_out0;
wire v_RD_7440_out0;
wire v_RD_7441_out0;
wire v_RD_7442_out0;
wire v_RD_7443_out0;
wire v_RD_7444_out0;
wire v_RD_7445_out0;
wire v_RD_7446_out0;
wire v_RD_7447_out0;
wire v_RD_7448_out0;
wire v_RD_7449_out0;
wire v_RD_7450_out0;
wire v_RD_7451_out0;
wire v_RD_7452_out0;
wire v_RD_7453_out0;
wire v_RD_7454_out0;
wire v_RD_7455_out0;
wire v_RD_7456_out0;
wire v_RD_7457_out0;
wire v_RD_7458_out0;
wire v_RD_7459_out0;
wire v_RD_7460_out0;
wire v_RD_7461_out0;
wire v_RD_7462_out0;
wire v_RD_7463_out0;
wire v_RD_7464_out0;
wire v_RD_7465_out0;
wire v_RD_7466_out0;
wire v_RD_7467_out0;
wire v_RD_7468_out0;
wire v_RD_7469_out0;
wire v_RD_7470_out0;
wire v_RD_7471_out0;
wire v_RD_7472_out0;
wire v_RD_7473_out0;
wire v_RD_7474_out0;
wire v_RD_7475_out0;
wire v_RD_7476_out0;
wire v_RD_7477_out0;
wire v_RD_7478_out0;
wire v_RD_7479_out0;
wire v_RD_7480_out0;
wire v_RD_7481_out0;
wire v_RD_7482_out0;
wire v_RD_7483_out0;
wire v_RD_7484_out0;
wire v_RD_7485_out0;
wire v_RD_7486_out0;
wire v_RD_7487_out0;
wire v_RD_7488_out0;
wire v_RD_7489_out0;
wire v_RD_7490_out0;
wire v_RD_7491_out0;
wire v_RD_7492_out0;
wire v_RD_7493_out0;
wire v_RD_7494_out0;
wire v_RD_7495_out0;
wire v_RD_7496_out0;
wire v_RD_7497_out0;
wire v_RD_7498_out0;
wire v_RD_7499_out0;
wire v_RD_7500_out0;
wire v_RD_7501_out0;
wire v_RD_7502_out0;
wire v_RD_7503_out0;
wire v_RD_7504_out0;
wire v_RD_7505_out0;
wire v_RD_7506_out0;
wire v_RD_7507_out0;
wire v_RD_7508_out0;
wire v_RD_7509_out0;
wire v_RD_7510_out0;
wire v_RD_7511_out0;
wire v_RD_7512_out0;
wire v_RD_7513_out0;
wire v_RD_7514_out0;
wire v_RD_7515_out0;
wire v_RD_7516_out0;
wire v_RD_7517_out0;
wire v_RD_7518_out0;
wire v_RD_7519_out0;
wire v_RD_7520_out0;
wire v_RD_7521_out0;
wire v_RD_7522_out0;
wire v_RD_7523_out0;
wire v_RD_7524_out0;
wire v_RD_7525_out0;
wire v_RD_7526_out0;
wire v_RD_7527_out0;
wire v_RD_7528_out0;
wire v_RD_7529_out0;
wire v_RD_7530_out0;
wire v_RD_7531_out0;
wire v_RD_7532_out0;
wire v_RD_7533_out0;
wire v_RD_7534_out0;
wire v_RD_7535_out0;
wire v_RD_7536_out0;
wire v_RD_7537_out0;
wire v_RD_7538_out0;
wire v_RD_7539_out0;
wire v_RD_7540_out0;
wire v_RD_7541_out0;
wire v_RD_7542_out0;
wire v_RD_7543_out0;
wire v_RD_7544_out0;
wire v_RD_7545_out0;
wire v_RD_7546_out0;
wire v_RD_7547_out0;
wire v_RD_7548_out0;
wire v_RD_7549_out0;
wire v_RD_7550_out0;
wire v_RD_7551_out0;
wire v_RD_7552_out0;
wire v_RD_7553_out0;
wire v_RD_7554_out0;
wire v_RD_7555_out0;
wire v_RD_7556_out0;
wire v_RD_7557_out0;
wire v_RD_7558_out0;
wire v_RD_7559_out0;
wire v_RD_7560_out0;
wire v_RD_7561_out0;
wire v_RD_7562_out0;
wire v_RD_7563_out0;
wire v_RD_7564_out0;
wire v_RD_7565_out0;
wire v_RD_7566_out0;
wire v_RD_7567_out0;
wire v_RD_7568_out0;
wire v_RD_7569_out0;
wire v_RD_7570_out0;
wire v_RD_7571_out0;
wire v_RD_7572_out0;
wire v_RD_7573_out0;
wire v_RD_7574_out0;
wire v_RD_7575_out0;
wire v_RD_7576_out0;
wire v_RD_7577_out0;
wire v_RD_7578_out0;
wire v_RD_7579_out0;
wire v_RD_7580_out0;
wire v_RD_7581_out0;
wire v_RD_7582_out0;
wire v_RD_7583_out0;
wire v_RD_7584_out0;
wire v_RD_7585_out0;
wire v_RD_7586_out0;
wire v_RD_7587_out0;
wire v_RD_7588_out0;
wire v_RD_7589_out0;
wire v_RD_7590_out0;
wire v_RD_7591_out0;
wire v_RD_7592_out0;
wire v_RD_7593_out0;
wire v_RD_7594_out0;
wire v_RD_7595_out0;
wire v_RD_7596_out0;
wire v_RD_7597_out0;
wire v_RD_7598_out0;
wire v_RD_7599_out0;
wire v_RD_7600_out0;
wire v_RD_7601_out0;
wire v_RD_7602_out0;
wire v_RD_7603_out0;
wire v_RD_7604_out0;
wire v_RD_7605_out0;
wire v_RD_7606_out0;
wire v_RD_7607_out0;
wire v_RD_7608_out0;
wire v_RD_7609_out0;
wire v_RD_7610_out0;
wire v_RD_7611_out0;
wire v_RD_7612_out0;
wire v_RD_7613_out0;
wire v_RD_7614_out0;
wire v_RD_7615_out0;
wire v_RD_7616_out0;
wire v_RD_7617_out0;
wire v_RD_7618_out0;
wire v_RD_7619_out0;
wire v_RD_7620_out0;
wire v_RD_7621_out0;
wire v_RD_7622_out0;
wire v_RD_7623_out0;
wire v_RD_7624_out0;
wire v_RD_7625_out0;
wire v_RD_7626_out0;
wire v_RD_7627_out0;
wire v_RD_7628_out0;
wire v_RD_7629_out0;
wire v_RD_7630_out0;
wire v_RD_7631_out0;
wire v_RD_7632_out0;
wire v_RD_7633_out0;
wire v_RD_7634_out0;
wire v_RD_SIGN_2405_out0;
wire v_RD_SIGN_2406_out0;
wire v_RD_SIGN_285_out0;
wire v_RD_SIGN_286_out0;
wire v_REN0_11136_out0;
wire v_REN1_6874_out0;
wire v_RESET_11174_out0;
wire v_RESET_11175_out0;
wire v_RESET_11176_out0;
wire v_RESET_11177_out0;
wire v_RESET_11178_out0;
wire v_RESET_11179_out0;
wire v_RESET_11180_out0;
wire v_RESET_11181_out0;
wire v_RESET_11182_out0;
wire v_RESET_11183_out0;
wire v_RESET_11184_out0;
wire v_RESET_11185_out0;
wire v_RESET_11186_out0;
wire v_RESET_11187_out0;
wire v_RESET_11188_out0;
wire v_RESET_11189_out0;
wire v_RM_11302_out0;
wire v_RM_11303_out0;
wire v_RM_11304_out0;
wire v_RM_11305_out0;
wire v_RM_11306_out0;
wire v_RM_11307_out0;
wire v_RM_11308_out0;
wire v_RM_11309_out0;
wire v_RM_11310_out0;
wire v_RM_11311_out0;
wire v_RM_11312_out0;
wire v_RM_11313_out0;
wire v_RM_11314_out0;
wire v_RM_11315_out0;
wire v_RM_11316_out0;
wire v_RM_11317_out0;
wire v_RM_11318_out0;
wire v_RM_11319_out0;
wire v_RM_11320_out0;
wire v_RM_11321_out0;
wire v_RM_11322_out0;
wire v_RM_11323_out0;
wire v_RM_11324_out0;
wire v_RM_11325_out0;
wire v_RM_11326_out0;
wire v_RM_11327_out0;
wire v_RM_11328_out0;
wire v_RM_11329_out0;
wire v_RM_11330_out0;
wire v_RM_11331_out0;
wire v_RM_11332_out0;
wire v_RM_11333_out0;
wire v_RM_11334_out0;
wire v_RM_11335_out0;
wire v_RM_11336_out0;
wire v_RM_11337_out0;
wire v_RM_11338_out0;
wire v_RM_11339_out0;
wire v_RM_11340_out0;
wire v_RM_11341_out0;
wire v_RM_11342_out0;
wire v_RM_11343_out0;
wire v_RM_11344_out0;
wire v_RM_11345_out0;
wire v_RM_11346_out0;
wire v_RM_11347_out0;
wire v_RM_11348_out0;
wire v_RM_11349_out0;
wire v_RM_11350_out0;
wire v_RM_11351_out0;
wire v_RM_11352_out0;
wire v_RM_11353_out0;
wire v_RM_11354_out0;
wire v_RM_11355_out0;
wire v_RM_11356_out0;
wire v_RM_11357_out0;
wire v_RM_11358_out0;
wire v_RM_11359_out0;
wire v_RM_11360_out0;
wire v_RM_11361_out0;
wire v_RM_11362_out0;
wire v_RM_11363_out0;
wire v_RM_11364_out0;
wire v_RM_11365_out0;
wire v_RM_11366_out0;
wire v_RM_11367_out0;
wire v_RM_11368_out0;
wire v_RM_11369_out0;
wire v_RM_11370_out0;
wire v_RM_11371_out0;
wire v_RM_11372_out0;
wire v_RM_11373_out0;
wire v_RM_11374_out0;
wire v_RM_11375_out0;
wire v_RM_11376_out0;
wire v_RM_11377_out0;
wire v_RM_11378_out0;
wire v_RM_11379_out0;
wire v_RM_11380_out0;
wire v_RM_11381_out0;
wire v_RM_11382_out0;
wire v_RM_11383_out0;
wire v_RM_11384_out0;
wire v_RM_11385_out0;
wire v_RM_11386_out0;
wire v_RM_11387_out0;
wire v_RM_11388_out0;
wire v_RM_11389_out0;
wire v_RM_11390_out0;
wire v_RM_11391_out0;
wire v_RM_11392_out0;
wire v_RM_11393_out0;
wire v_RM_11394_out0;
wire v_RM_11395_out0;
wire v_RM_11396_out0;
wire v_RM_11397_out0;
wire v_RM_11398_out0;
wire v_RM_11399_out0;
wire v_RM_11400_out0;
wire v_RM_11401_out0;
wire v_RM_11402_out0;
wire v_RM_11403_out0;
wire v_RM_11404_out0;
wire v_RM_11405_out0;
wire v_RM_11406_out0;
wire v_RM_11407_out0;
wire v_RM_11408_out0;
wire v_RM_11409_out0;
wire v_RM_11410_out0;
wire v_RM_11411_out0;
wire v_RM_11412_out0;
wire v_RM_11413_out0;
wire v_RM_11414_out0;
wire v_RM_11415_out0;
wire v_RM_11416_out0;
wire v_RM_11417_out0;
wire v_RM_11418_out0;
wire v_RM_11419_out0;
wire v_RM_11420_out0;
wire v_RM_11421_out0;
wire v_RM_11422_out0;
wire v_RM_11423_out0;
wire v_RM_11424_out0;
wire v_RM_11425_out0;
wire v_RM_11426_out0;
wire v_RM_11427_out0;
wire v_RM_11428_out0;
wire v_RM_11429_out0;
wire v_RM_11430_out0;
wire v_RM_11431_out0;
wire v_RM_11432_out0;
wire v_RM_11433_out0;
wire v_RM_11434_out0;
wire v_RM_11435_out0;
wire v_RM_11436_out0;
wire v_RM_11437_out0;
wire v_RM_11438_out0;
wire v_RM_11439_out0;
wire v_RM_11440_out0;
wire v_RM_11441_out0;
wire v_RM_11442_out0;
wire v_RM_11443_out0;
wire v_RM_11444_out0;
wire v_RM_11445_out0;
wire v_RM_11446_out0;
wire v_RM_11447_out0;
wire v_RM_11448_out0;
wire v_RM_11449_out0;
wire v_RM_11450_out0;
wire v_RM_11451_out0;
wire v_RM_11452_out0;
wire v_RM_11453_out0;
wire v_RM_11454_out0;
wire v_RM_11455_out0;
wire v_RM_11456_out0;
wire v_RM_11457_out0;
wire v_RM_11458_out0;
wire v_RM_11459_out0;
wire v_RM_11460_out0;
wire v_RM_11461_out0;
wire v_RM_11462_out0;
wire v_RM_11463_out0;
wire v_RM_11464_out0;
wire v_RM_11465_out0;
wire v_RM_11466_out0;
wire v_RM_11467_out0;
wire v_RM_11468_out0;
wire v_RM_11469_out0;
wire v_RM_11470_out0;
wire v_RM_11471_out0;
wire v_RM_11472_out0;
wire v_RM_11473_out0;
wire v_RM_11474_out0;
wire v_RM_11475_out0;
wire v_RM_11476_out0;
wire v_RM_11477_out0;
wire v_RM_11478_out0;
wire v_RM_11479_out0;
wire v_RM_11480_out0;
wire v_RM_11481_out0;
wire v_RM_11482_out0;
wire v_RM_11483_out0;
wire v_RM_11484_out0;
wire v_RM_11485_out0;
wire v_RM_11486_out0;
wire v_RM_11487_out0;
wire v_RM_11488_out0;
wire v_RM_11489_out0;
wire v_RM_11490_out0;
wire v_RM_11491_out0;
wire v_RM_11492_out0;
wire v_RM_11493_out0;
wire v_RM_11494_out0;
wire v_RM_11495_out0;
wire v_RM_11496_out0;
wire v_RM_11497_out0;
wire v_RM_11498_out0;
wire v_RM_11499_out0;
wire v_RM_11500_out0;
wire v_RM_11501_out0;
wire v_RM_11502_out0;
wire v_RM_11503_out0;
wire v_RM_11504_out0;
wire v_RM_11505_out0;
wire v_RM_11506_out0;
wire v_RM_11507_out0;
wire v_RM_11508_out0;
wire v_RM_11509_out0;
wire v_RM_11510_out0;
wire v_RM_11511_out0;
wire v_RM_11512_out0;
wire v_RM_11513_out0;
wire v_RM_11514_out0;
wire v_RM_11515_out0;
wire v_RM_11516_out0;
wire v_RM_11517_out0;
wire v_RM_11518_out0;
wire v_RM_11519_out0;
wire v_RM_11520_out0;
wire v_RM_11521_out0;
wire v_RM_11522_out0;
wire v_RM_11523_out0;
wire v_RM_11524_out0;
wire v_RM_11525_out0;
wire v_RM_11526_out0;
wire v_RM_11527_out0;
wire v_RM_11528_out0;
wire v_RM_11529_out0;
wire v_RM_11530_out0;
wire v_RM_11531_out0;
wire v_RM_11532_out0;
wire v_RM_11533_out0;
wire v_RM_11534_out0;
wire v_RM_11535_out0;
wire v_RM_11536_out0;
wire v_RM_11537_out0;
wire v_RM_11538_out0;
wire v_RM_11539_out0;
wire v_RM_11540_out0;
wire v_RM_11541_out0;
wire v_RM_11542_out0;
wire v_RM_11543_out0;
wire v_RM_11544_out0;
wire v_RM_11545_out0;
wire v_RM_11546_out0;
wire v_RM_11547_out0;
wire v_RM_11548_out0;
wire v_RM_11549_out0;
wire v_RM_11550_out0;
wire v_RM_11551_out0;
wire v_RM_11552_out0;
wire v_RM_11553_out0;
wire v_RM_11554_out0;
wire v_RM_11555_out0;
wire v_RM_11556_out0;
wire v_RM_11557_out0;
wire v_RM_11558_out0;
wire v_RM_11559_out0;
wire v_RM_11560_out0;
wire v_RM_11561_out0;
wire v_RM_11562_out0;
wire v_RM_11563_out0;
wire v_RM_11564_out0;
wire v_RM_11565_out0;
wire v_RM_11566_out0;
wire v_RM_11567_out0;
wire v_RM_11568_out0;
wire v_RM_11569_out0;
wire v_RM_11570_out0;
wire v_RM_11571_out0;
wire v_RM_11572_out0;
wire v_RM_11573_out0;
wire v_RM_11574_out0;
wire v_RM_11575_out0;
wire v_RM_11576_out0;
wire v_RM_11577_out0;
wire v_RM_11578_out0;
wire v_RM_11579_out0;
wire v_RM_11580_out0;
wire v_RM_11581_out0;
wire v_RM_11582_out0;
wire v_RM_11583_out0;
wire v_RM_11584_out0;
wire v_RM_11585_out0;
wire v_RM_11586_out0;
wire v_RM_11587_out0;
wire v_RM_11588_out0;
wire v_RM_11589_out0;
wire v_RM_11590_out0;
wire v_RM_11591_out0;
wire v_RM_11592_out0;
wire v_RM_11593_out0;
wire v_RM_11594_out0;
wire v_RM_11595_out0;
wire v_RM_11596_out0;
wire v_RM_11597_out0;
wire v_RM_11598_out0;
wire v_RM_11599_out0;
wire v_RM_11600_out0;
wire v_RM_11601_out0;
wire v_RM_11602_out0;
wire v_RM_11603_out0;
wire v_RM_11604_out0;
wire v_RM_11605_out0;
wire v_RM_11606_out0;
wire v_RM_11607_out0;
wire v_RM_11608_out0;
wire v_RM_11609_out0;
wire v_RM_11610_out0;
wire v_RM_11611_out0;
wire v_RM_11612_out0;
wire v_RM_11613_out0;
wire v_RM_11614_out0;
wire v_RM_11615_out0;
wire v_RM_11616_out0;
wire v_RM_11617_out0;
wire v_RM_11618_out0;
wire v_RM_11619_out0;
wire v_RM_11620_out0;
wire v_RM_11621_out0;
wire v_RM_11622_out0;
wire v_RM_11623_out0;
wire v_RM_11624_out0;
wire v_RM_11625_out0;
wire v_RM_11626_out0;
wire v_RM_11627_out0;
wire v_RM_11628_out0;
wire v_RM_11629_out0;
wire v_RM_11630_out0;
wire v_RM_11631_out0;
wire v_RM_11632_out0;
wire v_RM_11633_out0;
wire v_RM_11634_out0;
wire v_RM_11635_out0;
wire v_RM_11636_out0;
wire v_RM_11637_out0;
wire v_RM_11638_out0;
wire v_RM_11639_out0;
wire v_RM_11640_out0;
wire v_RM_11641_out0;
wire v_RM_11642_out0;
wire v_RM_11643_out0;
wire v_RM_11644_out0;
wire v_RM_11645_out0;
wire v_RM_11646_out0;
wire v_RM_11647_out0;
wire v_RM_11648_out0;
wire v_RM_11649_out0;
wire v_RM_11650_out0;
wire v_RM_11651_out0;
wire v_RM_11652_out0;
wire v_RM_11653_out0;
wire v_RM_11654_out0;
wire v_RM_11655_out0;
wire v_RM_11656_out0;
wire v_RM_11657_out0;
wire v_RM_11658_out0;
wire v_RM_11659_out0;
wire v_RM_11660_out0;
wire v_RM_11661_out0;
wire v_RM_11662_out0;
wire v_RM_11663_out0;
wire v_RM_11664_out0;
wire v_RM_11665_out0;
wire v_RM_11666_out0;
wire v_RM_11667_out0;
wire v_RM_11668_out0;
wire v_RM_11669_out0;
wire v_RM_11670_out0;
wire v_RM_11671_out0;
wire v_RM_11672_out0;
wire v_RM_11673_out0;
wire v_RM_11674_out0;
wire v_RM_11675_out0;
wire v_RM_11676_out0;
wire v_RM_11677_out0;
wire v_RM_11678_out0;
wire v_RM_11679_out0;
wire v_RM_11680_out0;
wire v_RM_11681_out0;
wire v_RM_11682_out0;
wire v_RM_11683_out0;
wire v_RM_11684_out0;
wire v_RM_11685_out0;
wire v_RM_11686_out0;
wire v_RM_11687_out0;
wire v_RM_11688_out0;
wire v_RM_11689_out0;
wire v_RM_11690_out0;
wire v_RM_11691_out0;
wire v_RM_11692_out0;
wire v_RM_11693_out0;
wire v_RM_11694_out0;
wire v_RM_11695_out0;
wire v_RM_11696_out0;
wire v_RM_11697_out0;
wire v_RM_11698_out0;
wire v_RM_11699_out0;
wire v_RM_11700_out0;
wire v_RM_11701_out0;
wire v_RM_11702_out0;
wire v_RM_11703_out0;
wire v_RM_11704_out0;
wire v_RM_11705_out0;
wire v_RM_11706_out0;
wire v_RM_11707_out0;
wire v_RM_11708_out0;
wire v_RM_11709_out0;
wire v_RM_11710_out0;
wire v_RM_11711_out0;
wire v_RM_11712_out0;
wire v_RM_11713_out0;
wire v_RM_11714_out0;
wire v_RM_11715_out0;
wire v_RM_11716_out0;
wire v_RM_11717_out0;
wire v_RM_11718_out0;
wire v_RM_11719_out0;
wire v_RM_11720_out0;
wire v_RM_11721_out0;
wire v_RM_11722_out0;
wire v_RM_11723_out0;
wire v_RM_11724_out0;
wire v_RM_11725_out0;
wire v_RM_11726_out0;
wire v_RM_11727_out0;
wire v_RM_11728_out0;
wire v_RM_11729_out0;
wire v_RM_11730_out0;
wire v_RM_11731_out0;
wire v_RM_11732_out0;
wire v_RM_11733_out0;
wire v_RM_11734_out0;
wire v_RM_11735_out0;
wire v_RM_11736_out0;
wire v_RM_11737_out0;
wire v_RM_11738_out0;
wire v_RM_11739_out0;
wire v_RM_11740_out0;
wire v_RM_11741_out0;
wire v_RM_11742_out0;
wire v_RM_11743_out0;
wire v_RM_11744_out0;
wire v_RM_11745_out0;
wire v_RM_11746_out0;
wire v_RM_11747_out0;
wire v_RM_11748_out0;
wire v_RM_11749_out0;
wire v_RM_11750_out0;
wire v_RM_11751_out0;
wire v_RM_11752_out0;
wire v_RM_11753_out0;
wire v_RM_11754_out0;
wire v_RM_11755_out0;
wire v_RM_11756_out0;
wire v_RM_11757_out0;
wire v_RM_11758_out0;
wire v_RM_11759_out0;
wire v_RM_11760_out0;
wire v_RM_11761_out0;
wire v_RM_11762_out0;
wire v_RM_11763_out0;
wire v_RM_11764_out0;
wire v_RM_11765_out0;
wire v_RM_11766_out0;
wire v_RM_11767_out0;
wire v_RM_11768_out0;
wire v_RM_11769_out0;
wire v_RM_11770_out0;
wire v_RM_11771_out0;
wire v_RM_11772_out0;
wire v_RM_11773_out0;
wire v_RM_11774_out0;
wire v_RM_11775_out0;
wire v_RM_11776_out0;
wire v_RM_11777_out0;
wire v_RM_11778_out0;
wire v_RM_11779_out0;
wire v_RM_11780_out0;
wire v_RM_11781_out0;
wire v_RM_11782_out0;
wire v_RM_11783_out0;
wire v_RM_11784_out0;
wire v_RM_11785_out0;
wire v_RM_11786_out0;
wire v_RM_11787_out0;
wire v_RM_11788_out0;
wire v_RM_11789_out0;
wire v_RM_11790_out0;
wire v_RM_11791_out0;
wire v_RM_11792_out0;
wire v_RM_11793_out0;
wire v_RM_11794_out0;
wire v_RM_11795_out0;
wire v_RM_11796_out0;
wire v_RM_11797_out0;
wire v_RM_11798_out0;
wire v_RM_11799_out0;
wire v_RM_11800_out0;
wire v_RM_11801_out0;
wire v_RM_11802_out0;
wire v_RM_11803_out0;
wire v_RM_11804_out0;
wire v_RM_11805_out0;
wire v_RM_11806_out0;
wire v_RM_11807_out0;
wire v_RM_11808_out0;
wire v_RM_11809_out0;
wire v_RM_11810_out0;
wire v_RM_11811_out0;
wire v_RM_11812_out0;
wire v_RM_11813_out0;
wire v_RM_11814_out0;
wire v_RM_11815_out0;
wire v_RM_11816_out0;
wire v_RM_11817_out0;
wire v_RM_11818_out0;
wire v_RM_11819_out0;
wire v_RM_11820_out0;
wire v_RM_11821_out0;
wire v_RM_11822_out0;
wire v_RM_11823_out0;
wire v_RM_11824_out0;
wire v_RM_11825_out0;
wire v_RM_11826_out0;
wire v_RM_11827_out0;
wire v_RM_11828_out0;
wire v_RM_11829_out0;
wire v_RM_11830_out0;
wire v_RM_11831_out0;
wire v_RM_11832_out0;
wire v_RM_11833_out0;
wire v_RM_11834_out0;
wire v_RM_11835_out0;
wire v_RM_11836_out0;
wire v_RM_11837_out0;
wire v_RM_11838_out0;
wire v_RM_11839_out0;
wire v_RM_11840_out0;
wire v_RM_11841_out0;
wire v_RM_11842_out0;
wire v_RM_11843_out0;
wire v_RM_11844_out0;
wire v_RM_11845_out0;
wire v_RM_11846_out0;
wire v_RM_11847_out0;
wire v_RM_11848_out0;
wire v_RM_11849_out0;
wire v_RM_11850_out0;
wire v_RM_11851_out0;
wire v_RM_11852_out0;
wire v_RM_11853_out0;
wire v_RM_11854_out0;
wire v_RM_11855_out0;
wire v_RM_11856_out0;
wire v_RM_11857_out0;
wire v_RM_11858_out0;
wire v_RM_11859_out0;
wire v_RM_11860_out0;
wire v_RM_11861_out0;
wire v_RM_11862_out0;
wire v_RM_11863_out0;
wire v_RM_11864_out0;
wire v_RM_11865_out0;
wire v_RM_11866_out0;
wire v_RM_11867_out0;
wire v_RM_11868_out0;
wire v_RM_11869_out0;
wire v_RM_11870_out0;
wire v_RM_11871_out0;
wire v_RM_11872_out0;
wire v_RM_11873_out0;
wire v_RM_11874_out0;
wire v_RM_11875_out0;
wire v_RM_11876_out0;
wire v_RM_11877_out0;
wire v_RM_11878_out0;
wire v_RM_11879_out0;
wire v_RM_11880_out0;
wire v_RM_11881_out0;
wire v_RM_11882_out0;
wire v_RM_11883_out0;
wire v_RM_11884_out0;
wire v_RM_11885_out0;
wire v_RM_11886_out0;
wire v_RM_11887_out0;
wire v_RM_11888_out0;
wire v_RM_11889_out0;
wire v_RM_11890_out0;
wire v_RM_11891_out0;
wire v_RM_11892_out0;
wire v_RM_11893_out0;
wire v_RM_11894_out0;
wire v_RM_11895_out0;
wire v_RM_11896_out0;
wire v_RM_11897_out0;
wire v_RM_11898_out0;
wire v_RM_11899_out0;
wire v_RM_11900_out0;
wire v_RM_11901_out0;
wire v_RM_11902_out0;
wire v_RM_11903_out0;
wire v_RM_11904_out0;
wire v_RM_11905_out0;
wire v_RM_11906_out0;
wire v_RM_11907_out0;
wire v_RM_11908_out0;
wire v_RM_11909_out0;
wire v_RM_11910_out0;
wire v_RM_11911_out0;
wire v_RM_11912_out0;
wire v_RM_11913_out0;
wire v_RM_11914_out0;
wire v_RM_11915_out0;
wire v_RM_11916_out0;
wire v_RM_11917_out0;
wire v_RM_11918_out0;
wire v_RM_11919_out0;
wire v_RM_11920_out0;
wire v_RM_11921_out0;
wire v_RM_11922_out0;
wire v_RM_11923_out0;
wire v_RM_11924_out0;
wire v_RM_11925_out0;
wire v_RM_11926_out0;
wire v_RM_11927_out0;
wire v_RM_11928_out0;
wire v_RM_11929_out0;
wire v_RM_11930_out0;
wire v_RM_11931_out0;
wire v_RM_11932_out0;
wire v_RM_11933_out0;
wire v_RM_11934_out0;
wire v_RM_11935_out0;
wire v_RM_11936_out0;
wire v_RM_11937_out0;
wire v_RM_11938_out0;
wire v_RM_11939_out0;
wire v_RM_11940_out0;
wire v_RM_11941_out0;
wire v_RM_11942_out0;
wire v_RM_11943_out0;
wire v_RM_11944_out0;
wire v_RM_11945_out0;
wire v_RM_11946_out0;
wire v_RM_11947_out0;
wire v_RM_11948_out0;
wire v_RM_11949_out0;
wire v_RM_11950_out0;
wire v_RM_11951_out0;
wire v_RM_11952_out0;
wire v_RM_11953_out0;
wire v_RM_11954_out0;
wire v_RM_11955_out0;
wire v_RM_11956_out0;
wire v_RM_11957_out0;
wire v_RM_11958_out0;
wire v_RM_11959_out0;
wire v_RM_11960_out0;
wire v_RM_11961_out0;
wire v_RM_11962_out0;
wire v_RM_11963_out0;
wire v_RM_11964_out0;
wire v_RM_11965_out0;
wire v_RM_11966_out0;
wire v_RM_11967_out0;
wire v_RM_11968_out0;
wire v_RM_11969_out0;
wire v_RM_11970_out0;
wire v_RM_11971_out0;
wire v_RM_11972_out0;
wire v_RM_11973_out0;
wire v_RM_11974_out0;
wire v_RM_11975_out0;
wire v_RM_11976_out0;
wire v_RM_11977_out0;
wire v_RM_11978_out0;
wire v_RM_11979_out0;
wire v_RM_11980_out0;
wire v_RM_11981_out0;
wire v_RM_11982_out0;
wire v_RM_11983_out0;
wire v_RM_11984_out0;
wire v_RM_11985_out0;
wire v_RM_11986_out0;
wire v_RM_11987_out0;
wire v_RM_11988_out0;
wire v_RM_11989_out0;
wire v_RM_11990_out0;
wire v_RM_11991_out0;
wire v_RM_11992_out0;
wire v_RM_11993_out0;
wire v_RM_11994_out0;
wire v_RM_11995_out0;
wire v_RM_11996_out0;
wire v_RM_11997_out0;
wire v_RM_11998_out0;
wire v_RM_11999_out0;
wire v_RM_12000_out0;
wire v_RM_12001_out0;
wire v_RM_12002_out0;
wire v_RM_12003_out0;
wire v_RM_12004_out0;
wire v_RM_12005_out0;
wire v_RM_12006_out0;
wire v_RM_12007_out0;
wire v_RM_12008_out0;
wire v_RM_12009_out0;
wire v_RM_12010_out0;
wire v_RM_12011_out0;
wire v_RM_12012_out0;
wire v_RM_12013_out0;
wire v_RM_12014_out0;
wire v_RM_12015_out0;
wire v_RM_12016_out0;
wire v_RM_12017_out0;
wire v_RM_12018_out0;
wire v_RM_12019_out0;
wire v_RM_12020_out0;
wire v_RM_12021_out0;
wire v_RM_12022_out0;
wire v_RM_12023_out0;
wire v_RM_12024_out0;
wire v_RM_12025_out0;
wire v_RM_12026_out0;
wire v_RM_12027_out0;
wire v_RM_12028_out0;
wire v_RM_12029_out0;
wire v_RM_12030_out0;
wire v_RM_12031_out0;
wire v_RM_12032_out0;
wire v_RM_12033_out0;
wire v_RM_12034_out0;
wire v_RM_12035_out0;
wire v_RM_12036_out0;
wire v_RM_12037_out0;
wire v_RM_12038_out0;
wire v_RM_12039_out0;
wire v_RM_12040_out0;
wire v_RM_12041_out0;
wire v_RM_12042_out0;
wire v_RM_12043_out0;
wire v_RM_12044_out0;
wire v_RM_12045_out0;
wire v_RM_12046_out0;
wire v_RM_12047_out0;
wire v_RM_12048_out0;
wire v_RM_12049_out0;
wire v_RM_12050_out0;
wire v_RM_12051_out0;
wire v_RM_12052_out0;
wire v_RM_12053_out0;
wire v_RM_12054_out0;
wire v_RM_12055_out0;
wire v_RM_12056_out0;
wire v_RM_12057_out0;
wire v_RM_12058_out0;
wire v_RM_12059_out0;
wire v_RM_12060_out0;
wire v_RM_12061_out0;
wire v_RM_12062_out0;
wire v_RM_12063_out0;
wire v_RM_12064_out0;
wire v_RM_12065_out0;
wire v_RM_12066_out0;
wire v_RM_12067_out0;
wire v_RM_12068_out0;
wire v_RM_12069_out0;
wire v_RM_12070_out0;
wire v_RM_12071_out0;
wire v_RM_12072_out0;
wire v_RM_12073_out0;
wire v_RM_12074_out0;
wire v_RM_12075_out0;
wire v_RM_12076_out0;
wire v_RM_12077_out0;
wire v_RM_12078_out0;
wire v_RM_12079_out0;
wire v_RM_12080_out0;
wire v_RM_12081_out0;
wire v_RM_12082_out0;
wire v_RM_12083_out0;
wire v_RM_12084_out0;
wire v_RM_12085_out0;
wire v_RM_12086_out0;
wire v_RM_12087_out0;
wire v_RM_12088_out0;
wire v_RM_12089_out0;
wire v_RM_12090_out0;
wire v_RM_12091_out0;
wire v_RM_12092_out0;
wire v_RM_12093_out0;
wire v_RM_12094_out0;
wire v_RM_12095_out0;
wire v_RM_12096_out0;
wire v_RM_12097_out0;
wire v_RM_12098_out0;
wire v_RM_12099_out0;
wire v_RM_12100_out0;
wire v_RM_12101_out0;
wire v_RM_12102_out0;
wire v_RM_12103_out0;
wire v_RM_12104_out0;
wire v_RM_12105_out0;
wire v_RM_12106_out0;
wire v_RM_12107_out0;
wire v_RM_12108_out0;
wire v_RM_12109_out0;
wire v_RM_12110_out0;
wire v_RM_12111_out0;
wire v_RM_12112_out0;
wire v_RM_12113_out0;
wire v_RM_12114_out0;
wire v_RM_12115_out0;
wire v_RM_12116_out0;
wire v_RM_12117_out0;
wire v_RM_12118_out0;
wire v_RM_12119_out0;
wire v_RM_12120_out0;
wire v_RM_12121_out0;
wire v_RM_12122_out0;
wire v_RM_12123_out0;
wire v_RM_12124_out0;
wire v_RM_12125_out0;
wire v_RM_12126_out0;
wire v_RM_12127_out0;
wire v_RM_12128_out0;
wire v_RM_12129_out0;
wire v_RM_12130_out0;
wire v_RM_12131_out0;
wire v_RM_12132_out0;
wire v_RM_12133_out0;
wire v_RM_12134_out0;
wire v_RM_12135_out0;
wire v_RM_12136_out0;
wire v_RM_12137_out0;
wire v_RM_12138_out0;
wire v_RM_12139_out0;
wire v_RM_12140_out0;
wire v_RM_12141_out0;
wire v_RM_12142_out0;
wire v_RM_12143_out0;
wire v_RM_12144_out0;
wire v_RM_12145_out0;
wire v_RM_12146_out0;
wire v_RM_12147_out0;
wire v_RM_12148_out0;
wire v_RM_12149_out0;
wire v_RM_12150_out0;
wire v_RM_12151_out0;
wire v_RM_12152_out0;
wire v_RM_12153_out0;
wire v_RM_12154_out0;
wire v_RM_12155_out0;
wire v_RM_12156_out0;
wire v_RM_12157_out0;
wire v_RM_12158_out0;
wire v_RM_12159_out0;
wire v_RM_12160_out0;
wire v_RM_12161_out0;
wire v_RM_12162_out0;
wire v_RM_12163_out0;
wire v_RM_12164_out0;
wire v_RM_12165_out0;
wire v_RM_12166_out0;
wire v_RM_12167_out0;
wire v_RM_12168_out0;
wire v_RM_12169_out0;
wire v_RM_12170_out0;
wire v_RM_12171_out0;
wire v_RM_12172_out0;
wire v_RM_12173_out0;
wire v_RM_12174_out0;
wire v_RM_12175_out0;
wire v_RM_12176_out0;
wire v_RM_12177_out0;
wire v_RM_12178_out0;
wire v_RM_12179_out0;
wire v_RM_12180_out0;
wire v_RM_12181_out0;
wire v_RM_12182_out0;
wire v_RM_12183_out0;
wire v_RM_12184_out0;
wire v_RM_12185_out0;
wire v_RM_12186_out0;
wire v_RM_12187_out0;
wire v_RM_12188_out0;
wire v_RM_12189_out0;
wire v_RM_12190_out0;
wire v_RM_12191_out0;
wire v_RM_12192_out0;
wire v_RM_12193_out0;
wire v_RM_12194_out0;
wire v_RM_12195_out0;
wire v_RM_12196_out0;
wire v_RM_12197_out0;
wire v_RM_12198_out0;
wire v_RM_12199_out0;
wire v_RM_12200_out0;
wire v_RM_12201_out0;
wire v_RM_12202_out0;
wire v_RM_12203_out0;
wire v_RM_12204_out0;
wire v_RM_12205_out0;
wire v_RM_12206_out0;
wire v_RM_12207_out0;
wire v_RM_12208_out0;
wire v_RM_12209_out0;
wire v_RM_12210_out0;
wire v_RM_12211_out0;
wire v_RM_12212_out0;
wire v_RM_12213_out0;
wire v_RM_12214_out0;
wire v_RM_12215_out0;
wire v_RM_12216_out0;
wire v_RM_12217_out0;
wire v_RM_12218_out0;
wire v_RM_12219_out0;
wire v_RM_12220_out0;
wire v_RM_12221_out0;
wire v_RM_12222_out0;
wire v_RM_12223_out0;
wire v_RM_12224_out0;
wire v_RM_12225_out0;
wire v_RM_12226_out0;
wire v_RM_12227_out0;
wire v_RM_12228_out0;
wire v_RM_12229_out0;
wire v_RM_3355_out0;
wire v_RM_3356_out0;
wire v_RM_3357_out0;
wire v_RM_3358_out0;
wire v_RM_3359_out0;
wire v_RM_3360_out0;
wire v_RM_3361_out0;
wire v_RM_3362_out0;
wire v_RM_3363_out0;
wire v_RM_3364_out0;
wire v_RM_3365_out0;
wire v_RM_3366_out0;
wire v_RM_3367_out0;
wire v_RM_3368_out0;
wire v_RM_3369_out0;
wire v_RM_3370_out0;
wire v_RM_3371_out0;
wire v_RM_3372_out0;
wire v_RM_3373_out0;
wire v_RM_3374_out0;
wire v_RM_3375_out0;
wire v_RM_3376_out0;
wire v_RM_3377_out0;
wire v_RM_3378_out0;
wire v_RM_3379_out0;
wire v_RM_3380_out0;
wire v_RM_3381_out0;
wire v_RM_3382_out0;
wire v_RM_3383_out0;
wire v_RM_3384_out0;
wire v_RM_3385_out0;
wire v_RM_3386_out0;
wire v_RM_3387_out0;
wire v_RM_3388_out0;
wire v_RM_3389_out0;
wire v_RM_3390_out0;
wire v_RM_3391_out0;
wire v_RM_3392_out0;
wire v_RM_3393_out0;
wire v_RM_3394_out0;
wire v_RM_3395_out0;
wire v_RM_3396_out0;
wire v_RM_3397_out0;
wire v_RM_3398_out0;
wire v_RM_3399_out0;
wire v_RM_3400_out0;
wire v_RM_3401_out0;
wire v_RM_3402_out0;
wire v_RM_3403_out0;
wire v_RM_3404_out0;
wire v_RM_3405_out0;
wire v_RM_3406_out0;
wire v_RM_3407_out0;
wire v_RM_3408_out0;
wire v_RM_3409_out0;
wire v_RM_3410_out0;
wire v_RM_3411_out0;
wire v_RM_3412_out0;
wire v_RM_3413_out0;
wire v_RM_3414_out0;
wire v_RM_3415_out0;
wire v_RM_3416_out0;
wire v_RM_3417_out0;
wire v_RM_3418_out0;
wire v_RM_3419_out0;
wire v_RM_3420_out0;
wire v_RM_3421_out0;
wire v_RM_3422_out0;
wire v_RM_3423_out0;
wire v_RM_3424_out0;
wire v_RM_3425_out0;
wire v_RM_3426_out0;
wire v_RM_3427_out0;
wire v_RM_3428_out0;
wire v_RM_3429_out0;
wire v_RM_3430_out0;
wire v_RM_3431_out0;
wire v_RM_3432_out0;
wire v_RM_3433_out0;
wire v_RM_3434_out0;
wire v_RM_3435_out0;
wire v_RM_3436_out0;
wire v_RM_3437_out0;
wire v_RM_3438_out0;
wire v_RM_3439_out0;
wire v_RM_3440_out0;
wire v_RM_3441_out0;
wire v_RM_3442_out0;
wire v_RM_3443_out0;
wire v_RM_3444_out0;
wire v_RM_3445_out0;
wire v_RM_3446_out0;
wire v_RM_3447_out0;
wire v_RM_3448_out0;
wire v_RM_3449_out0;
wire v_RM_3450_out0;
wire v_RM_3451_out0;
wire v_RM_3452_out0;
wire v_RM_3453_out0;
wire v_RM_3454_out0;
wire v_RM_3455_out0;
wire v_RM_3456_out0;
wire v_RM_3457_out0;
wire v_RM_3458_out0;
wire v_RM_3459_out0;
wire v_RM_3460_out0;
wire v_RM_3461_out0;
wire v_RM_3462_out0;
wire v_RM_3463_out0;
wire v_RM_3464_out0;
wire v_RM_3465_out0;
wire v_RM_3466_out0;
wire v_RM_3467_out0;
wire v_RM_3468_out0;
wire v_RM_3469_out0;
wire v_RM_3470_out0;
wire v_RM_3471_out0;
wire v_RM_3472_out0;
wire v_RM_3473_out0;
wire v_RM_3474_out0;
wire v_RM_3475_out0;
wire v_RM_3476_out0;
wire v_RM_3477_out0;
wire v_RM_3478_out0;
wire v_RM_3479_out0;
wire v_RM_3480_out0;
wire v_RM_3481_out0;
wire v_RM_3482_out0;
wire v_RM_3483_out0;
wire v_RM_3484_out0;
wire v_RM_3485_out0;
wire v_RM_3486_out0;
wire v_RM_3487_out0;
wire v_RM_3488_out0;
wire v_RM_3489_out0;
wire v_RM_3490_out0;
wire v_RM_3491_out0;
wire v_RM_3492_out0;
wire v_RM_3493_out0;
wire v_RM_3494_out0;
wire v_RM_3495_out0;
wire v_RM_3496_out0;
wire v_RM_3497_out0;
wire v_RM_3498_out0;
wire v_RM_3499_out0;
wire v_RM_3500_out0;
wire v_RM_3501_out0;
wire v_RM_3502_out0;
wire v_RM_3503_out0;
wire v_RM_3504_out0;
wire v_RM_3505_out0;
wire v_RM_3506_out0;
wire v_RM_3507_out0;
wire v_RM_3508_out0;
wire v_RM_3509_out0;
wire v_RM_3510_out0;
wire v_RM_3511_out0;
wire v_RM_3512_out0;
wire v_RM_3513_out0;
wire v_RM_3514_out0;
wire v_RM_3515_out0;
wire v_RM_3516_out0;
wire v_RM_3517_out0;
wire v_RM_3518_out0;
wire v_RM_3519_out0;
wire v_RM_3520_out0;
wire v_RM_3521_out0;
wire v_RM_3522_out0;
wire v_RM_3523_out0;
wire v_RM_3524_out0;
wire v_RM_3525_out0;
wire v_RM_3526_out0;
wire v_RM_3527_out0;
wire v_RM_3528_out0;
wire v_RM_3529_out0;
wire v_RM_3530_out0;
wire v_RM_3531_out0;
wire v_RM_3532_out0;
wire v_RM_3533_out0;
wire v_RM_3534_out0;
wire v_RM_3535_out0;
wire v_RM_3536_out0;
wire v_RM_3537_out0;
wire v_RM_3538_out0;
wire v_RM_3539_out0;
wire v_RM_3540_out0;
wire v_RM_3541_out0;
wire v_RM_3542_out0;
wire v_RM_3543_out0;
wire v_RM_3544_out0;
wire v_RM_3545_out0;
wire v_RM_3546_out0;
wire v_RM_3547_out0;
wire v_RM_3548_out0;
wire v_RM_3549_out0;
wire v_RM_3550_out0;
wire v_RM_3551_out0;
wire v_RM_3552_out0;
wire v_RM_3553_out0;
wire v_RM_3554_out0;
wire v_RM_3555_out0;
wire v_RM_3556_out0;
wire v_RM_3557_out0;
wire v_RM_3558_out0;
wire v_RM_3559_out0;
wire v_RM_3560_out0;
wire v_RM_3561_out0;
wire v_RM_3562_out0;
wire v_RM_3563_out0;
wire v_RM_3564_out0;
wire v_RM_3565_out0;
wire v_RM_3566_out0;
wire v_RM_3567_out0;
wire v_RM_3568_out0;
wire v_RM_3569_out0;
wire v_RM_3570_out0;
wire v_RM_3571_out0;
wire v_RM_3572_out0;
wire v_RM_3573_out0;
wire v_RM_3574_out0;
wire v_RM_3575_out0;
wire v_RM_3576_out0;
wire v_RM_3577_out0;
wire v_RM_3578_out0;
wire v_RM_3579_out0;
wire v_RM_3580_out0;
wire v_RM_3581_out0;
wire v_RM_3582_out0;
wire v_RM_3583_out0;
wire v_RM_3584_out0;
wire v_RM_3585_out0;
wire v_RM_3586_out0;
wire v_RM_3587_out0;
wire v_RM_3588_out0;
wire v_RM_3589_out0;
wire v_RM_3590_out0;
wire v_RM_3591_out0;
wire v_RM_3592_out0;
wire v_RM_3593_out0;
wire v_RM_3594_out0;
wire v_RM_3595_out0;
wire v_RM_3596_out0;
wire v_RM_3597_out0;
wire v_RM_3598_out0;
wire v_RM_3599_out0;
wire v_RM_3600_out0;
wire v_RM_3601_out0;
wire v_RM_3602_out0;
wire v_RM_3603_out0;
wire v_RM_3604_out0;
wire v_RM_3605_out0;
wire v_RM_3606_out0;
wire v_RM_3607_out0;
wire v_RM_3608_out0;
wire v_RM_3609_out0;
wire v_RM_3610_out0;
wire v_RM_3611_out0;
wire v_RM_3612_out0;
wire v_RM_3613_out0;
wire v_RM_3614_out0;
wire v_RM_3615_out0;
wire v_RM_3616_out0;
wire v_RM_3617_out0;
wire v_RM_3618_out0;
wire v_RM_3619_out0;
wire v_RM_3620_out0;
wire v_RM_3621_out0;
wire v_RM_3622_out0;
wire v_RM_3623_out0;
wire v_RM_3624_out0;
wire v_RM_3625_out0;
wire v_RM_3626_out0;
wire v_RM_3627_out0;
wire v_RM_3628_out0;
wire v_RM_3629_out0;
wire v_RM_3630_out0;
wire v_RM_3631_out0;
wire v_RM_3632_out0;
wire v_RM_3633_out0;
wire v_RM_3634_out0;
wire v_RM_3635_out0;
wire v_RM_3636_out0;
wire v_RM_3637_out0;
wire v_RM_3638_out0;
wire v_RM_3639_out0;
wire v_RM_3640_out0;
wire v_RM_3641_out0;
wire v_RM_3642_out0;
wire v_RM_3643_out0;
wire v_RM_3644_out0;
wire v_RM_3645_out0;
wire v_RM_3646_out0;
wire v_RM_3647_out0;
wire v_RM_3648_out0;
wire v_RM_3649_out0;
wire v_RM_3650_out0;
wire v_RM_3651_out0;
wire v_RM_3652_out0;
wire v_RM_3653_out0;
wire v_RM_3654_out0;
wire v_RM_3655_out0;
wire v_RM_3656_out0;
wire v_RM_3657_out0;
wire v_RM_3658_out0;
wire v_RM_3659_out0;
wire v_RM_3660_out0;
wire v_RM_3661_out0;
wire v_RM_3662_out0;
wire v_RM_3663_out0;
wire v_RM_3664_out0;
wire v_RM_3665_out0;
wire v_RM_3666_out0;
wire v_RM_3667_out0;
wire v_RM_3668_out0;
wire v_RM_3669_out0;
wire v_RM_3670_out0;
wire v_RM_3671_out0;
wire v_RM_3672_out0;
wire v_RM_3673_out0;
wire v_RM_3674_out0;
wire v_RM_3675_out0;
wire v_RM_3676_out0;
wire v_RM_3677_out0;
wire v_RM_3678_out0;
wire v_RM_3679_out0;
wire v_RM_3680_out0;
wire v_RM_3681_out0;
wire v_RM_3682_out0;
wire v_RM_3683_out0;
wire v_RM_3684_out0;
wire v_RM_3685_out0;
wire v_RM_3686_out0;
wire v_RM_3687_out0;
wire v_RM_3688_out0;
wire v_RM_3689_out0;
wire v_RM_3690_out0;
wire v_RM_3691_out0;
wire v_RM_3692_out0;
wire v_RM_3693_out0;
wire v_RM_3694_out0;
wire v_RM_3695_out0;
wire v_RM_3696_out0;
wire v_RM_3697_out0;
wire v_RM_3698_out0;
wire v_RM_3699_out0;
wire v_RM_3700_out0;
wire v_RM_3701_out0;
wire v_RM_3702_out0;
wire v_RM_3703_out0;
wire v_RM_3704_out0;
wire v_RM_3705_out0;
wire v_RM_3706_out0;
wire v_RM_3707_out0;
wire v_RM_3708_out0;
wire v_RM_3709_out0;
wire v_RM_3710_out0;
wire v_RM_3711_out0;
wire v_RM_3712_out0;
wire v_RM_3713_out0;
wire v_RM_3714_out0;
wire v_RM_3715_out0;
wire v_RM_3716_out0;
wire v_RM_3717_out0;
wire v_RM_3718_out0;
wire v_RM_3719_out0;
wire v_RM_3720_out0;
wire v_RM_3721_out0;
wire v_RM_3722_out0;
wire v_RM_3723_out0;
wire v_RM_3724_out0;
wire v_RM_3725_out0;
wire v_RM_3726_out0;
wire v_RM_3727_out0;
wire v_RM_3728_out0;
wire v_RM_3729_out0;
wire v_RM_3730_out0;
wire v_RM_3731_out0;
wire v_RM_3732_out0;
wire v_RM_3733_out0;
wire v_RM_3734_out0;
wire v_RM_3735_out0;
wire v_RM_3736_out0;
wire v_RM_3737_out0;
wire v_RM_3738_out0;
wire v_RM_3739_out0;
wire v_RM_3740_out0;
wire v_RM_3741_out0;
wire v_RM_3742_out0;
wire v_RM_3743_out0;
wire v_RM_3744_out0;
wire v_RM_3745_out0;
wire v_RM_3746_out0;
wire v_RM_3747_out0;
wire v_RM_3748_out0;
wire v_RM_3749_out0;
wire v_RM_3750_out0;
wire v_RM_3751_out0;
wire v_RM_3752_out0;
wire v_RM_3753_out0;
wire v_RM_3754_out0;
wire v_RM_3755_out0;
wire v_RM_3756_out0;
wire v_RM_3757_out0;
wire v_RM_3758_out0;
wire v_RM_3759_out0;
wire v_RM_3760_out0;
wire v_RM_3761_out0;
wire v_RM_3762_out0;
wire v_RM_3763_out0;
wire v_RM_3764_out0;
wire v_RM_3765_out0;
wire v_RM_3766_out0;
wire v_RM_3767_out0;
wire v_RM_3768_out0;
wire v_RM_3769_out0;
wire v_RM_3770_out0;
wire v_RM_3771_out0;
wire v_RM_3772_out0;
wire v_RM_3773_out0;
wire v_RM_3774_out0;
wire v_RM_3775_out0;
wire v_RM_3776_out0;
wire v_RM_3777_out0;
wire v_RM_3778_out0;
wire v_RM_3779_out0;
wire v_RM_3780_out0;
wire v_RM_3781_out0;
wire v_RM_3782_out0;
wire v_RM_3783_out0;
wire v_RM_3784_out0;
wire v_RM_3785_out0;
wire v_RM_3786_out0;
wire v_RM_3787_out0;
wire v_RM_3788_out0;
wire v_RM_3789_out0;
wire v_RM_3790_out0;
wire v_RM_3791_out0;
wire v_RM_3792_out0;
wire v_RM_3793_out0;
wire v_RM_3794_out0;
wire v_RM_3795_out0;
wire v_RM_3796_out0;
wire v_RM_3797_out0;
wire v_RM_3798_out0;
wire v_RM_3799_out0;
wire v_RM_3800_out0;
wire v_RM_3801_out0;
wire v_RM_3802_out0;
wire v_ROM1_462_out0;
wire v_ROR_282_out0;
wire v_ROR_283_out0;
wire v_ROR_3286_out0;
wire v_ROR_3287_out0;
wire v_ROR_3288_out0;
wire v_ROR_3289_out0;
wire v_ROR_544_out0;
wire v_ROR_545_out0;
wire v_RXBYTERECEIVED_3269_out0;
wire v_RXBYTERECEIVED_91_out0;
wire v_RX_BYTEREADY_8756_out0;
wire v_RX_BYTE_READY_2436_out0;
wire v_RX_DONE_RECEIVING_10484_out0;
wire v_RX_INST0_2970_out0;
wire v_RX_INST1_12_out0;
wire v_RX_INSTRUCTION_11170_out0;
wire v_RX_INSTRUCTION_11171_out0;
wire v_RX_INSTRUCTION_13325_out0;
wire v_RX_INSTRUCTION_2343_out0;
wire v_RX_INSTRUCTION_2344_out0;
wire v_RX_INSTRUCTION_3258_out0;
wire v_RX_INSTRUCTION_3259_out0;
wire v_RX_INSTRUCTION_4659_out0;
wire v_RX_INSTRUCTION_8686_out0;
wire v_RX_INSTRUCTION_94_out0;
wire v_RX_INSTRUCTION_95_out0;
wire v_RX_INST_2334_out0;
wire v_RX_OVERFLOW_426_out0;
wire v_RX_OVERFLOW_4469_out0;
wire v_RX_OVERFLOW_5848_out0;
wire v_SBC_11051_out0;
wire v_SBC_11052_out0;
wire v_SBC_13605_out0;
wire v_SBC_13606_out0;
wire v_SBC_4825_out0;
wire v_SBC_4826_out0;
wire v_SEL1_10304_out0;
wire v_SEL1_1164_out0;
wire v_SEL1_1204_out0;
wire v_SEL1_13445_out0;
wire v_SEL1_2305_out0;
wire v_SEL1_2306_out0;
wire v_SEL1_2319_out0;
wire v_SEL1_240_out0;
wire v_SEL1_2428_out0;
wire v_SEL1_2914_out0;
wire v_SEL1_2915_out0;
wire v_SEL1_4858_out0;
wire v_SEL2_10323_out0;
wire v_SEL2_10324_out0;
wire v_SEL2_280_out0;
wire v_SEL2_281_out0;
wire v_SEL3_1143_out0;
wire v_SEL3_1144_out0;
wire v_SEL3_2615_out0;
wire v_SEL3_2616_out0;
wire v_SEL4_7636_out0;
wire v_SEL4_7637_out0;
wire v_SEL5_3049_out0;
wire v_SEL5_3050_out0;
wire v_SHIFHT_ENABLE_13500_out0;
wire v_SHIFHT_ENABLE_13501_out0;
wire v_SHIFHT_ENABLE_13502_out0;
wire v_SHIFHT_ENABLE_13503_out0;
wire v_SHIFT_ENABLE_8684_out0;
wire v_SHIFT_RD_2544_out0;
wire v_SHIFT_RD_2545_out0;
wire v_SHIFT_WHICH_OP_10465_out0;
wire v_SHIFT_WHICH_OP_10466_out0;
wire v_SHIFT_WHICH_OP_10715_out0;
wire v_SHIFT_WHICH_OP_10716_out0;
wire v_SHIFT_WHICH_OP_4459_out0;
wire v_SHIFT_WHICH_OP_4460_out0;
wire v_SIGN_ANS_10302_out0;
wire v_SIGN_ANS_10303_out0;
wire v_SIGN_ANS_1970_out0;
wire v_SIGN_ANS_1971_out0;
wire v_SIGN_ANS_4457_out0;
wire v_SIGN_ANS_4458_out0;
wire v_SIGN_ANS_8650_out0;
wire v_SIGN_ANS_8651_out0;
wire v_STALL_10281_out0;
wire v_STALL_10282_out0;
wire v_STALL_1758_out0;
wire v_STALL_1759_out0;
wire v_STALL_427_out0;
wire v_STALL_428_out0;
wire v_STALL_6910_out0;
wire v_STALL_6911_out0;
wire v_STALL_DUAL_CORE_12234_out0;
wire v_STALL_DUAL_CORE_12235_out0;
wire v_STALL_DUAL_CORE_13617_out0;
wire v_STALL_DUAL_CORE_13618_out0;
wire v_STALL_DUAL_CORE_1738_out0;
wire v_STALL_DUAL_CORE_1739_out0;
wire v_STALL_DUAL_CORE_1958_out0;
wire v_STALL_DUAL_CORE_1959_out0;
wire v_STALL_DUAL_CORE_3127_out0;
wire v_STALL_DUAL_CORE_3128_out0;
wire v_STALL_DUAL_CORE_3264_out0;
wire v_STALL_DUAL_CORE_3265_out0;
wire v_STALL_DUAL_CORE_4695_out0;
wire v_STALL_DUAL_CORE_4696_out0;
wire v_STALL_dual_core_8741_out0;
wire v_STALL_dual_core_8742_out0;
wire v_STARTBIT_6967_out0;
wire v_STARTBIT_6968_out0;
wire v_STARTBIT_6969_out0;
wire v_STARTBIT_6970_out0;
wire v_START_13394_out0;
wire v_START_13395_out0;
wire v_START_3027_out0;
wire v_START_3028_out0;
wire v_START_392_out0;
wire v_START_393_out0;
wire v_STAT_INSTRUCTION_10272_out0;
wire v_STAT_INSTRUCTION_10273_out0;
wire v_STAT_INSTRUCTION_2434_out0;
wire v_STAT_INSTRUCTION_2435_out0;
wire v_STAT_INSTRUCTION_2855_out0;
wire v_STAT_INSTRUCTION_2856_out0;
wire v_STORE_10831_out0;
wire v_STORE_10832_out0;
wire v_STORE_1195_out0;
wire v_STORE_1196_out0;
wire v_STORE_12245_out0;
wire v_STORE_12246_out0;
wire v_STORE_13298_out0;
wire v_STORE_13299_out0;
wire v_STORE_221_out0;
wire v_STORE_222_out0;
wire v_STORE_540_out0;
wire v_STORE_541_out0;
wire v_STORE_PCOUNTER_2102_out0;
wire v_STORE_PCOUNTER_2103_out0;
wire v_STORE_WEN_4544_out0;
wire v_STORE_WEN_4545_out0;
wire v_STORE_pccounter_2883_out0;
wire v_STORE_pccounter_2884_out0;
wire v_STP_10307_out0;
wire v_STP_10308_out0;
wire v_STP_10352_out0;
wire v_STP_10353_out0;
wire v_STP_10467_out0;
wire v_STP_10468_out0;
wire v_STP_10977_out0;
wire v_STP_10978_out0;
wire v_STP_11240_out0;
wire v_STP_11241_out0;
wire v_STP_52_out0;
wire v_STP_53_out0;
wire v_SUBNORMAL_8808_out0;
wire v_SUBNORMAL_8809_out0;
wire v_SUB_12247_out0;
wire v_SUB_12248_out0;
wire v_SUB_2695_out0;
wire v_SUB_2696_out0;
wire v_SUB_2909_out0;
wire v_SUB_2910_out0;
wire v_SUB_2957_out0;
wire v_SUB_2958_out0;
wire v_SUB_4616_out0;
wire v_SUB_4617_out0;
wire v_SUB_4618_out0;
wire v_SUB_4619_out0;
wire v_SUB_8663_out0;
wire v_SUB_8664_out0;
wire v_SUB_INSTRUCTION_11195_out0;
wire v_SUB_INSTRUCTION_11196_out0;
wire v_SUB_INSTRUCTION_2789_out0;
wire v_SUB_INSTRUCTION_2790_out0;
wire v_SUB_INSTRUCTION_7085_out0;
wire v_SUB_INSTRUCTION_7086_out0;
wire v_S_11300_out0;
wire v_S_11301_out0;
wire v_S_1219_out0;
wire v_S_1220_out0;
wire v_S_1221_out0;
wire v_S_1222_out0;
wire v_S_1223_out0;
wire v_S_1224_out0;
wire v_S_1225_out0;
wire v_S_1226_out0;
wire v_S_1227_out0;
wire v_S_1228_out0;
wire v_S_1229_out0;
wire v_S_1230_out0;
wire v_S_1231_out0;
wire v_S_1232_out0;
wire v_S_1233_out0;
wire v_S_1234_out0;
wire v_S_1235_out0;
wire v_S_1236_out0;
wire v_S_1237_out0;
wire v_S_1238_out0;
wire v_S_1239_out0;
wire v_S_1240_out0;
wire v_S_1241_out0;
wire v_S_1242_out0;
wire v_S_1243_out0;
wire v_S_1244_out0;
wire v_S_1245_out0;
wire v_S_1246_out0;
wire v_S_1247_out0;
wire v_S_1248_out0;
wire v_S_1249_out0;
wire v_S_1250_out0;
wire v_S_1251_out0;
wire v_S_1252_out0;
wire v_S_1253_out0;
wire v_S_1254_out0;
wire v_S_1255_out0;
wire v_S_1256_out0;
wire v_S_1257_out0;
wire v_S_1258_out0;
wire v_S_1259_out0;
wire v_S_1260_out0;
wire v_S_1261_out0;
wire v_S_1262_out0;
wire v_S_1263_out0;
wire v_S_1264_out0;
wire v_S_1265_out0;
wire v_S_1266_out0;
wire v_S_1267_out0;
wire v_S_1268_out0;
wire v_S_1269_out0;
wire v_S_1270_out0;
wire v_S_1271_out0;
wire v_S_1272_out0;
wire v_S_1273_out0;
wire v_S_1274_out0;
wire v_S_1275_out0;
wire v_S_1276_out0;
wire v_S_1277_out0;
wire v_S_1278_out0;
wire v_S_1279_out0;
wire v_S_1280_out0;
wire v_S_1281_out0;
wire v_S_1282_out0;
wire v_S_1283_out0;
wire v_S_1284_out0;
wire v_S_1285_out0;
wire v_S_1286_out0;
wire v_S_1287_out0;
wire v_S_1288_out0;
wire v_S_1289_out0;
wire v_S_1290_out0;
wire v_S_1291_out0;
wire v_S_1292_out0;
wire v_S_1293_out0;
wire v_S_1294_out0;
wire v_S_1295_out0;
wire v_S_1296_out0;
wire v_S_1297_out0;
wire v_S_1298_out0;
wire v_S_1299_out0;
wire v_S_1300_out0;
wire v_S_1301_out0;
wire v_S_1302_out0;
wire v_S_1303_out0;
wire v_S_1304_out0;
wire v_S_1305_out0;
wire v_S_1306_out0;
wire v_S_1307_out0;
wire v_S_1308_out0;
wire v_S_1309_out0;
wire v_S_1310_out0;
wire v_S_1311_out0;
wire v_S_1312_out0;
wire v_S_1313_out0;
wire v_S_1314_out0;
wire v_S_1315_out0;
wire v_S_1316_out0;
wire v_S_1317_out0;
wire v_S_1318_out0;
wire v_S_1319_out0;
wire v_S_1320_out0;
wire v_S_1321_out0;
wire v_S_1322_out0;
wire v_S_1323_out0;
wire v_S_1324_out0;
wire v_S_1325_out0;
wire v_S_1326_out0;
wire v_S_1327_out0;
wire v_S_1328_out0;
wire v_S_1329_out0;
wire v_S_1330_out0;
wire v_S_1331_out0;
wire v_S_1332_out0;
wire v_S_1333_out0;
wire v_S_1334_out0;
wire v_S_1335_out0;
wire v_S_1336_out0;
wire v_S_1337_out0;
wire v_S_1338_out0;
wire v_S_1339_out0;
wire v_S_1340_out0;
wire v_S_1341_out0;
wire v_S_1342_out0;
wire v_S_1343_out0;
wire v_S_1344_out0;
wire v_S_1345_out0;
wire v_S_1346_out0;
wire v_S_1347_out0;
wire v_S_1348_out0;
wire v_S_1349_out0;
wire v_S_1350_out0;
wire v_S_1351_out0;
wire v_S_1352_out0;
wire v_S_1353_out0;
wire v_S_1354_out0;
wire v_S_1355_out0;
wire v_S_1356_out0;
wire v_S_1357_out0;
wire v_S_1358_out0;
wire v_S_1359_out0;
wire v_S_1360_out0;
wire v_S_1361_out0;
wire v_S_1362_out0;
wire v_S_1363_out0;
wire v_S_1364_out0;
wire v_S_1365_out0;
wire v_S_1366_out0;
wire v_S_1367_out0;
wire v_S_1368_out0;
wire v_S_1369_out0;
wire v_S_1370_out0;
wire v_S_1371_out0;
wire v_S_1372_out0;
wire v_S_1373_out0;
wire v_S_1374_out0;
wire v_S_1375_out0;
wire v_S_1376_out0;
wire v_S_1377_out0;
wire v_S_1378_out0;
wire v_S_1379_out0;
wire v_S_1380_out0;
wire v_S_1381_out0;
wire v_S_1382_out0;
wire v_S_1383_out0;
wire v_S_1384_out0;
wire v_S_1385_out0;
wire v_S_1386_out0;
wire v_S_1387_out0;
wire v_S_1388_out0;
wire v_S_1389_out0;
wire v_S_1390_out0;
wire v_S_1391_out0;
wire v_S_1392_out0;
wire v_S_1393_out0;
wire v_S_1394_out0;
wire v_S_1395_out0;
wire v_S_1396_out0;
wire v_S_1397_out0;
wire v_S_1398_out0;
wire v_S_1399_out0;
wire v_S_1400_out0;
wire v_S_1401_out0;
wire v_S_1402_out0;
wire v_S_1403_out0;
wire v_S_1404_out0;
wire v_S_1405_out0;
wire v_S_1406_out0;
wire v_S_1407_out0;
wire v_S_1408_out0;
wire v_S_1409_out0;
wire v_S_1410_out0;
wire v_S_1411_out0;
wire v_S_1412_out0;
wire v_S_1413_out0;
wire v_S_1414_out0;
wire v_S_1415_out0;
wire v_S_1416_out0;
wire v_S_1417_out0;
wire v_S_1418_out0;
wire v_S_1419_out0;
wire v_S_1420_out0;
wire v_S_1421_out0;
wire v_S_1422_out0;
wire v_S_1423_out0;
wire v_S_1424_out0;
wire v_S_1425_out0;
wire v_S_1426_out0;
wire v_S_1427_out0;
wire v_S_1428_out0;
wire v_S_1429_out0;
wire v_S_1430_out0;
wire v_S_1431_out0;
wire v_S_1432_out0;
wire v_S_1433_out0;
wire v_S_1434_out0;
wire v_S_1435_out0;
wire v_S_1436_out0;
wire v_S_1437_out0;
wire v_S_1438_out0;
wire v_S_1439_out0;
wire v_S_1440_out0;
wire v_S_1441_out0;
wire v_S_1442_out0;
wire v_S_1443_out0;
wire v_S_1444_out0;
wire v_S_1445_out0;
wire v_S_1446_out0;
wire v_S_1447_out0;
wire v_S_1448_out0;
wire v_S_1449_out0;
wire v_S_1450_out0;
wire v_S_1451_out0;
wire v_S_1452_out0;
wire v_S_1453_out0;
wire v_S_1454_out0;
wire v_S_1455_out0;
wire v_S_1456_out0;
wire v_S_1457_out0;
wire v_S_1458_out0;
wire v_S_1459_out0;
wire v_S_1460_out0;
wire v_S_1461_out0;
wire v_S_1462_out0;
wire v_S_1463_out0;
wire v_S_1464_out0;
wire v_S_1465_out0;
wire v_S_1466_out0;
wire v_S_1467_out0;
wire v_S_1468_out0;
wire v_S_1469_out0;
wire v_S_1470_out0;
wire v_S_1471_out0;
wire v_S_1472_out0;
wire v_S_1473_out0;
wire v_S_1474_out0;
wire v_S_1475_out0;
wire v_S_1476_out0;
wire v_S_1477_out0;
wire v_S_1478_out0;
wire v_S_1479_out0;
wire v_S_1480_out0;
wire v_S_1481_out0;
wire v_S_1482_out0;
wire v_S_1483_out0;
wire v_S_1484_out0;
wire v_S_1485_out0;
wire v_S_1486_out0;
wire v_S_1487_out0;
wire v_S_1488_out0;
wire v_S_1489_out0;
wire v_S_1490_out0;
wire v_S_1491_out0;
wire v_S_1492_out0;
wire v_S_1493_out0;
wire v_S_1494_out0;
wire v_S_1495_out0;
wire v_S_1496_out0;
wire v_S_1497_out0;
wire v_S_1498_out0;
wire v_S_1499_out0;
wire v_S_1500_out0;
wire v_S_1501_out0;
wire v_S_1502_out0;
wire v_S_1503_out0;
wire v_S_1504_out0;
wire v_S_1505_out0;
wire v_S_1506_out0;
wire v_S_1507_out0;
wire v_S_1508_out0;
wire v_S_1509_out0;
wire v_S_1510_out0;
wire v_S_1511_out0;
wire v_S_1512_out0;
wire v_S_1513_out0;
wire v_S_1514_out0;
wire v_S_1515_out0;
wire v_S_1516_out0;
wire v_S_1517_out0;
wire v_S_1518_out0;
wire v_S_1519_out0;
wire v_S_1520_out0;
wire v_S_1521_out0;
wire v_S_1522_out0;
wire v_S_1523_out0;
wire v_S_1524_out0;
wire v_S_1525_out0;
wire v_S_1526_out0;
wire v_S_1527_out0;
wire v_S_1528_out0;
wire v_S_1529_out0;
wire v_S_1530_out0;
wire v_S_1531_out0;
wire v_S_1532_out0;
wire v_S_1533_out0;
wire v_S_1534_out0;
wire v_S_1535_out0;
wire v_S_1536_out0;
wire v_S_1537_out0;
wire v_S_1538_out0;
wire v_S_1539_out0;
wire v_S_1540_out0;
wire v_S_1541_out0;
wire v_S_1542_out0;
wire v_S_1543_out0;
wire v_S_1544_out0;
wire v_S_1545_out0;
wire v_S_1546_out0;
wire v_S_1547_out0;
wire v_S_1548_out0;
wire v_S_1549_out0;
wire v_S_1550_out0;
wire v_S_1551_out0;
wire v_S_1552_out0;
wire v_S_1553_out0;
wire v_S_1554_out0;
wire v_S_1555_out0;
wire v_S_1556_out0;
wire v_S_1557_out0;
wire v_S_1558_out0;
wire v_S_1559_out0;
wire v_S_1560_out0;
wire v_S_1561_out0;
wire v_S_1562_out0;
wire v_S_1563_out0;
wire v_S_1564_out0;
wire v_S_1565_out0;
wire v_S_1566_out0;
wire v_S_1567_out0;
wire v_S_1568_out0;
wire v_S_1569_out0;
wire v_S_1570_out0;
wire v_S_1571_out0;
wire v_S_1572_out0;
wire v_S_1573_out0;
wire v_S_1574_out0;
wire v_S_1575_out0;
wire v_S_1576_out0;
wire v_S_1577_out0;
wire v_S_1578_out0;
wire v_S_1579_out0;
wire v_S_1580_out0;
wire v_S_1581_out0;
wire v_S_1582_out0;
wire v_S_1583_out0;
wire v_S_1584_out0;
wire v_S_1585_out0;
wire v_S_1586_out0;
wire v_S_1587_out0;
wire v_S_1588_out0;
wire v_S_1589_out0;
wire v_S_1590_out0;
wire v_S_1591_out0;
wire v_S_1592_out0;
wire v_S_1593_out0;
wire v_S_1594_out0;
wire v_S_1595_out0;
wire v_S_1596_out0;
wire v_S_1597_out0;
wire v_S_1598_out0;
wire v_S_1599_out0;
wire v_S_1600_out0;
wire v_S_1601_out0;
wire v_S_1602_out0;
wire v_S_1603_out0;
wire v_S_1604_out0;
wire v_S_1605_out0;
wire v_S_1606_out0;
wire v_S_1607_out0;
wire v_S_1608_out0;
wire v_S_1609_out0;
wire v_S_1610_out0;
wire v_S_1611_out0;
wire v_S_1612_out0;
wire v_S_1613_out0;
wire v_S_1614_out0;
wire v_S_1615_out0;
wire v_S_1616_out0;
wire v_S_1617_out0;
wire v_S_1618_out0;
wire v_S_1619_out0;
wire v_S_1620_out0;
wire v_S_1621_out0;
wire v_S_1622_out0;
wire v_S_1623_out0;
wire v_S_1624_out0;
wire v_S_1625_out0;
wire v_S_1626_out0;
wire v_S_1627_out0;
wire v_S_1628_out0;
wire v_S_1629_out0;
wire v_S_1630_out0;
wire v_S_1631_out0;
wire v_S_1632_out0;
wire v_S_1633_out0;
wire v_S_1634_out0;
wire v_S_1635_out0;
wire v_S_1636_out0;
wire v_S_1637_out0;
wire v_S_1638_out0;
wire v_S_1639_out0;
wire v_S_1640_out0;
wire v_S_1641_out0;
wire v_S_1642_out0;
wire v_S_1643_out0;
wire v_S_1644_out0;
wire v_S_1645_out0;
wire v_S_1646_out0;
wire v_S_1647_out0;
wire v_S_1648_out0;
wire v_S_1649_out0;
wire v_S_1650_out0;
wire v_S_1651_out0;
wire v_S_1652_out0;
wire v_S_1653_out0;
wire v_S_1654_out0;
wire v_S_1655_out0;
wire v_S_1656_out0;
wire v_S_1657_out0;
wire v_S_1658_out0;
wire v_S_1659_out0;
wire v_S_1660_out0;
wire v_S_1661_out0;
wire v_S_1662_out0;
wire v_S_1663_out0;
wire v_S_1664_out0;
wire v_S_1665_out0;
wire v_S_1666_out0;
wire v_S_4665_out0;
wire v_S_4666_out0;
wire v_S_4667_out0;
wire v_S_4668_out0;
wire v_S_4669_out0;
wire v_S_4670_out0;
wire v_S_4671_out0;
wire v_S_4672_out0;
wire v_S_4673_out0;
wire v_S_4674_out0;
wire v_S_4675_out0;
wire v_S_4676_out0;
wire v_S_4677_out0;
wire v_S_4678_out0;
wire v_S_4679_out0;
wire v_S_4680_out0;
wire v_S_4681_out0;
wire v_S_4682_out0;
wire v_S_4683_out0;
wire v_S_4684_out0;
wire v_S_4685_out0;
wire v_S_4686_out0;
wire v_S_4687_out0;
wire v_S_4688_out0;
wire v_S_4689_out0;
wire v_S_4690_out0;
wire v_S_4691_out0;
wire v_S_4692_out0;
wire v_S_4693_out0;
wire v_S_4694_out0;
wire v_S_8863_out0;
wire v_S_8864_out0;
wire v_S_8865_out0;
wire v_S_8866_out0;
wire v_S_8867_out0;
wire v_S_8868_out0;
wire v_S_8869_out0;
wire v_S_8870_out0;
wire v_S_8871_out0;
wire v_S_8872_out0;
wire v_S_8873_out0;
wire v_S_8874_out0;
wire v_S_8875_out0;
wire v_S_8876_out0;
wire v_S_8877_out0;
wire v_S_8878_out0;
wire v_S_8879_out0;
wire v_S_8880_out0;
wire v_S_8881_out0;
wire v_S_8882_out0;
wire v_S_8883_out0;
wire v_S_8884_out0;
wire v_S_8885_out0;
wire v_S_8886_out0;
wire v_S_8887_out0;
wire v_S_8888_out0;
wire v_S_8889_out0;
wire v_S_8890_out0;
wire v_S_8891_out0;
wire v_S_8892_out0;
wire v_S_8893_out0;
wire v_S_8894_out0;
wire v_S_8895_out0;
wire v_S_8896_out0;
wire v_S_8897_out0;
wire v_S_8898_out0;
wire v_S_8899_out0;
wire v_S_8900_out0;
wire v_S_8901_out0;
wire v_S_8902_out0;
wire v_S_8903_out0;
wire v_S_8904_out0;
wire v_S_8905_out0;
wire v_S_8906_out0;
wire v_S_8907_out0;
wire v_S_8908_out0;
wire v_S_8909_out0;
wire v_S_8910_out0;
wire v_S_8911_out0;
wire v_S_8912_out0;
wire v_S_8913_out0;
wire v_S_8914_out0;
wire v_S_8915_out0;
wire v_S_8916_out0;
wire v_S_8917_out0;
wire v_S_8918_out0;
wire v_S_8919_out0;
wire v_S_8920_out0;
wire v_S_8921_out0;
wire v_S_8922_out0;
wire v_S_8923_out0;
wire v_S_8924_out0;
wire v_S_8925_out0;
wire v_S_8926_out0;
wire v_S_8927_out0;
wire v_S_8928_out0;
wire v_S_8929_out0;
wire v_S_8930_out0;
wire v_S_8931_out0;
wire v_S_8932_out0;
wire v_S_8933_out0;
wire v_S_8934_out0;
wire v_S_8935_out0;
wire v_S_8936_out0;
wire v_S_8937_out0;
wire v_S_8938_out0;
wire v_S_8939_out0;
wire v_S_8940_out0;
wire v_S_8941_out0;
wire v_S_8942_out0;
wire v_S_8943_out0;
wire v_S_8944_out0;
wire v_S_8945_out0;
wire v_S_8946_out0;
wire v_S_8947_out0;
wire v_S_8948_out0;
wire v_S_8949_out0;
wire v_S_8950_out0;
wire v_S_8951_out0;
wire v_S_8952_out0;
wire v_S_8953_out0;
wire v_S_8954_out0;
wire v_S_8955_out0;
wire v_S_8956_out0;
wire v_S_8957_out0;
wire v_S_8958_out0;
wire v_S_8959_out0;
wire v_S_8960_out0;
wire v_S_8961_out0;
wire v_S_8962_out0;
wire v_S_8963_out0;
wire v_S_8964_out0;
wire v_S_8965_out0;
wire v_S_8966_out0;
wire v_S_8967_out0;
wire v_S_8968_out0;
wire v_S_8969_out0;
wire v_S_8970_out0;
wire v_S_8971_out0;
wire v_S_8972_out0;
wire v_S_8973_out0;
wire v_S_8974_out0;
wire v_S_8975_out0;
wire v_S_8976_out0;
wire v_S_8977_out0;
wire v_S_8978_out0;
wire v_S_8979_out0;
wire v_S_8980_out0;
wire v_S_8981_out0;
wire v_S_8982_out0;
wire v_S_8983_out0;
wire v_S_8984_out0;
wire v_S_8985_out0;
wire v_S_8986_out0;
wire v_S_8987_out0;
wire v_S_8988_out0;
wire v_S_8989_out0;
wire v_S_8990_out0;
wire v_S_8991_out0;
wire v_S_8992_out0;
wire v_S_8993_out0;
wire v_S_8994_out0;
wire v_S_8995_out0;
wire v_S_8996_out0;
wire v_S_8997_out0;
wire v_S_8998_out0;
wire v_S_8999_out0;
wire v_S_9000_out0;
wire v_S_9001_out0;
wire v_S_9002_out0;
wire v_S_9003_out0;
wire v_S_9004_out0;
wire v_S_9005_out0;
wire v_S_9006_out0;
wire v_S_9007_out0;
wire v_S_9008_out0;
wire v_S_9009_out0;
wire v_S_9010_out0;
wire v_S_9011_out0;
wire v_S_9012_out0;
wire v_S_9013_out0;
wire v_S_9014_out0;
wire v_S_9015_out0;
wire v_S_9016_out0;
wire v_S_9017_out0;
wire v_S_9018_out0;
wire v_S_9019_out0;
wire v_S_9020_out0;
wire v_S_9021_out0;
wire v_S_9022_out0;
wire v_S_9023_out0;
wire v_S_9024_out0;
wire v_S_9025_out0;
wire v_S_9026_out0;
wire v_S_9027_out0;
wire v_S_9028_out0;
wire v_S_9029_out0;
wire v_S_9030_out0;
wire v_S_9031_out0;
wire v_S_9032_out0;
wire v_S_9033_out0;
wire v_S_9034_out0;
wire v_S_9035_out0;
wire v_S_9036_out0;
wire v_S_9037_out0;
wire v_S_9038_out0;
wire v_S_9039_out0;
wire v_S_9040_out0;
wire v_S_9041_out0;
wire v_S_9042_out0;
wire v_S_9043_out0;
wire v_S_9044_out0;
wire v_S_9045_out0;
wire v_S_9046_out0;
wire v_S_9047_out0;
wire v_S_9048_out0;
wire v_S_9049_out0;
wire v_S_9050_out0;
wire v_S_9051_out0;
wire v_S_9052_out0;
wire v_S_9053_out0;
wire v_S_9054_out0;
wire v_S_9055_out0;
wire v_S_9056_out0;
wire v_S_9057_out0;
wire v_S_9058_out0;
wire v_S_9059_out0;
wire v_S_9060_out0;
wire v_S_9061_out0;
wire v_S_9062_out0;
wire v_S_9063_out0;
wire v_S_9064_out0;
wire v_S_9065_out0;
wire v_S_9066_out0;
wire v_S_9067_out0;
wire v_S_9068_out0;
wire v_S_9069_out0;
wire v_S_9070_out0;
wire v_S_9071_out0;
wire v_S_9072_out0;
wire v_S_9073_out0;
wire v_S_9074_out0;
wire v_S_9075_out0;
wire v_S_9076_out0;
wire v_S_9077_out0;
wire v_S_9078_out0;
wire v_S_9079_out0;
wire v_S_9080_out0;
wire v_S_9081_out0;
wire v_S_9082_out0;
wire v_S_9083_out0;
wire v_S_9084_out0;
wire v_S_9085_out0;
wire v_S_9086_out0;
wire v_S_9087_out0;
wire v_S_9088_out0;
wire v_S_9089_out0;
wire v_S_9090_out0;
wire v_S_9091_out0;
wire v_S_9092_out0;
wire v_S_9093_out0;
wire v_S_9094_out0;
wire v_S_9095_out0;
wire v_S_9096_out0;
wire v_S_9097_out0;
wire v_S_9098_out0;
wire v_S_9099_out0;
wire v_S_9100_out0;
wire v_S_9101_out0;
wire v_S_9102_out0;
wire v_S_9103_out0;
wire v_S_9104_out0;
wire v_S_9105_out0;
wire v_S_9106_out0;
wire v_S_9107_out0;
wire v_S_9108_out0;
wire v_S_9109_out0;
wire v_S_9110_out0;
wire v_S_9111_out0;
wire v_S_9112_out0;
wire v_S_9113_out0;
wire v_S_9114_out0;
wire v_S_9115_out0;
wire v_S_9116_out0;
wire v_S_9117_out0;
wire v_S_9118_out0;
wire v_S_9119_out0;
wire v_S_9120_out0;
wire v_S_9121_out0;
wire v_S_9122_out0;
wire v_S_9123_out0;
wire v_S_9124_out0;
wire v_S_9125_out0;
wire v_S_9126_out0;
wire v_S_9127_out0;
wire v_S_9128_out0;
wire v_S_9129_out0;
wire v_S_9130_out0;
wire v_S_9131_out0;
wire v_S_9132_out0;
wire v_S_9133_out0;
wire v_S_9134_out0;
wire v_S_9135_out0;
wire v_S_9136_out0;
wire v_S_9137_out0;
wire v_S_9138_out0;
wire v_S_9139_out0;
wire v_S_9140_out0;
wire v_S_9141_out0;
wire v_S_9142_out0;
wire v_S_9143_out0;
wire v_S_9144_out0;
wire v_S_9145_out0;
wire v_S_9146_out0;
wire v_S_9147_out0;
wire v_S_9148_out0;
wire v_S_9149_out0;
wire v_S_9150_out0;
wire v_S_9151_out0;
wire v_S_9152_out0;
wire v_S_9153_out0;
wire v_S_9154_out0;
wire v_S_9155_out0;
wire v_S_9156_out0;
wire v_S_9157_out0;
wire v_S_9158_out0;
wire v_S_9159_out0;
wire v_S_9160_out0;
wire v_S_9161_out0;
wire v_S_9162_out0;
wire v_S_9163_out0;
wire v_S_9164_out0;
wire v_S_9165_out0;
wire v_S_9166_out0;
wire v_S_9167_out0;
wire v_S_9168_out0;
wire v_S_9169_out0;
wire v_S_9170_out0;
wire v_S_9171_out0;
wire v_S_9172_out0;
wire v_S_9173_out0;
wire v_S_9174_out0;
wire v_S_9175_out0;
wire v_S_9176_out0;
wire v_S_9177_out0;
wire v_S_9178_out0;
wire v_S_9179_out0;
wire v_S_9180_out0;
wire v_S_9181_out0;
wire v_S_9182_out0;
wire v_S_9183_out0;
wire v_S_9184_out0;
wire v_S_9185_out0;
wire v_S_9186_out0;
wire v_S_9187_out0;
wire v_S_9188_out0;
wire v_S_9189_out0;
wire v_S_9190_out0;
wire v_S_9191_out0;
wire v_S_9192_out0;
wire v_S_9193_out0;
wire v_S_9194_out0;
wire v_S_9195_out0;
wire v_S_9196_out0;
wire v_S_9197_out0;
wire v_S_9198_out0;
wire v_S_9199_out0;
wire v_S_9200_out0;
wire v_S_9201_out0;
wire v_S_9202_out0;
wire v_S_9203_out0;
wire v_S_9204_out0;
wire v_S_9205_out0;
wire v_S_9206_out0;
wire v_S_9207_out0;
wire v_S_9208_out0;
wire v_S_9209_out0;
wire v_S_9210_out0;
wire v_S_9211_out0;
wire v_S_9212_out0;
wire v_S_9213_out0;
wire v_S_9214_out0;
wire v_S_9215_out0;
wire v_S_9216_out0;
wire v_S_9217_out0;
wire v_S_9218_out0;
wire v_S_9219_out0;
wire v_S_9220_out0;
wire v_S_9221_out0;
wire v_S_9222_out0;
wire v_S_9223_out0;
wire v_S_9224_out0;
wire v_S_9225_out0;
wire v_S_9226_out0;
wire v_S_9227_out0;
wire v_S_9228_out0;
wire v_S_9229_out0;
wire v_S_9230_out0;
wire v_S_9231_out0;
wire v_S_9232_out0;
wire v_S_9233_out0;
wire v_S_9234_out0;
wire v_S_9235_out0;
wire v_S_9236_out0;
wire v_S_9237_out0;
wire v_S_9238_out0;
wire v_S_9239_out0;
wire v_S_9240_out0;
wire v_S_9241_out0;
wire v_S_9242_out0;
wire v_S_9243_out0;
wire v_S_9244_out0;
wire v_S_9245_out0;
wire v_S_9246_out0;
wire v_S_9247_out0;
wire v_S_9248_out0;
wire v_S_9249_out0;
wire v_S_9250_out0;
wire v_S_9251_out0;
wire v_S_9252_out0;
wire v_S_9253_out0;
wire v_S_9254_out0;
wire v_S_9255_out0;
wire v_S_9256_out0;
wire v_S_9257_out0;
wire v_S_9258_out0;
wire v_S_9259_out0;
wire v_S_9260_out0;
wire v_S_9261_out0;
wire v_S_9262_out0;
wire v_S_9263_out0;
wire v_S_9264_out0;
wire v_S_9265_out0;
wire v_S_9266_out0;
wire v_S_9267_out0;
wire v_S_9268_out0;
wire v_S_9269_out0;
wire v_S_9270_out0;
wire v_S_9271_out0;
wire v_S_9272_out0;
wire v_S_9273_out0;
wire v_S_9274_out0;
wire v_S_9275_out0;
wire v_S_9276_out0;
wire v_S_9277_out0;
wire v_S_9278_out0;
wire v_S_9279_out0;
wire v_S_9280_out0;
wire v_S_9281_out0;
wire v_S_9282_out0;
wire v_S_9283_out0;
wire v_S_9284_out0;
wire v_S_9285_out0;
wire v_S_9286_out0;
wire v_S_9287_out0;
wire v_S_9288_out0;
wire v_S_9289_out0;
wire v_S_9290_out0;
wire v_S_9291_out0;
wire v_S_9292_out0;
wire v_S_9293_out0;
wire v_S_9294_out0;
wire v_S_9295_out0;
wire v_S_9296_out0;
wire v_S_9297_out0;
wire v_S_9298_out0;
wire v_S_9299_out0;
wire v_S_9300_out0;
wire v_S_9301_out0;
wire v_S_9302_out0;
wire v_S_9303_out0;
wire v_S_9304_out0;
wire v_S_9305_out0;
wire v_S_9306_out0;
wire v_S_9307_out0;
wire v_S_9308_out0;
wire v_S_9309_out0;
wire v_S_9310_out0;
wire v_S_9311_out0;
wire v_S_9312_out0;
wire v_S_9313_out0;
wire v_S_9314_out0;
wire v_S_9315_out0;
wire v_S_9316_out0;
wire v_S_9317_out0;
wire v_S_9318_out0;
wire v_S_9319_out0;
wire v_S_9320_out0;
wire v_S_9321_out0;
wire v_S_9322_out0;
wire v_S_9323_out0;
wire v_S_9324_out0;
wire v_S_9325_out0;
wire v_S_9326_out0;
wire v_S_9327_out0;
wire v_S_9328_out0;
wire v_S_9329_out0;
wire v_S_9330_out0;
wire v_S_9331_out0;
wire v_S_9332_out0;
wire v_S_9333_out0;
wire v_S_9334_out0;
wire v_S_9335_out0;
wire v_S_9336_out0;
wire v_S_9337_out0;
wire v_S_9338_out0;
wire v_S_9339_out0;
wire v_S_9340_out0;
wire v_S_9341_out0;
wire v_S_9342_out0;
wire v_S_9343_out0;
wire v_S_9344_out0;
wire v_S_9345_out0;
wire v_S_9346_out0;
wire v_S_9347_out0;
wire v_S_9348_out0;
wire v_S_9349_out0;
wire v_S_9350_out0;
wire v_S_9351_out0;
wire v_S_9352_out0;
wire v_S_9353_out0;
wire v_S_9354_out0;
wire v_S_9355_out0;
wire v_S_9356_out0;
wire v_S_9357_out0;
wire v_S_9358_out0;
wire v_S_9359_out0;
wire v_S_9360_out0;
wire v_S_9361_out0;
wire v_S_9362_out0;
wire v_S_9363_out0;
wire v_S_9364_out0;
wire v_S_9365_out0;
wire v_S_9366_out0;
wire v_S_9367_out0;
wire v_S_9368_out0;
wire v_S_9369_out0;
wire v_S_9370_out0;
wire v_S_9371_out0;
wire v_S_9372_out0;
wire v_S_9373_out0;
wire v_S_9374_out0;
wire v_S_9375_out0;
wire v_S_9376_out0;
wire v_S_9377_out0;
wire v_S_9378_out0;
wire v_S_9379_out0;
wire v_S_9380_out0;
wire v_S_9381_out0;
wire v_S_9382_out0;
wire v_S_9383_out0;
wire v_S_9384_out0;
wire v_S_9385_out0;
wire v_S_9386_out0;
wire v_S_9387_out0;
wire v_S_9388_out0;
wire v_S_9389_out0;
wire v_S_9390_out0;
wire v_S_9391_out0;
wire v_S_9392_out0;
wire v_S_9393_out0;
wire v_S_9394_out0;
wire v_S_9395_out0;
wire v_S_9396_out0;
wire v_S_9397_out0;
wire v_S_9398_out0;
wire v_S_9399_out0;
wire v_S_9400_out0;
wire v_S_9401_out0;
wire v_S_9402_out0;
wire v_S_9403_out0;
wire v_S_9404_out0;
wire v_S_9405_out0;
wire v_S_9406_out0;
wire v_S_9407_out0;
wire v_S_9408_out0;
wire v_S_9409_out0;
wire v_S_9410_out0;
wire v_S_9411_out0;
wire v_S_9412_out0;
wire v_S_9413_out0;
wire v_S_9414_out0;
wire v_S_9415_out0;
wire v_S_9416_out0;
wire v_S_9417_out0;
wire v_S_9418_out0;
wire v_S_9419_out0;
wire v_S_9420_out0;
wire v_S_9421_out0;
wire v_S_9422_out0;
wire v_S_9423_out0;
wire v_S_9424_out0;
wire v_S_9425_out0;
wire v_S_9426_out0;
wire v_S_9427_out0;
wire v_S_9428_out0;
wire v_S_9429_out0;
wire v_S_9430_out0;
wire v_S_9431_out0;
wire v_S_9432_out0;
wire v_S_9433_out0;
wire v_S_9434_out0;
wire v_S_9435_out0;
wire v_S_9436_out0;
wire v_S_9437_out0;
wire v_S_9438_out0;
wire v_S_9439_out0;
wire v_S_9440_out0;
wire v_S_9441_out0;
wire v_S_9442_out0;
wire v_S_9443_out0;
wire v_S_9444_out0;
wire v_S_9445_out0;
wire v_S_9446_out0;
wire v_S_9447_out0;
wire v_S_9448_out0;
wire v_S_9449_out0;
wire v_S_9450_out0;
wire v_S_9451_out0;
wire v_S_9452_out0;
wire v_S_9453_out0;
wire v_S_9454_out0;
wire v_S_9455_out0;
wire v_S_9456_out0;
wire v_S_9457_out0;
wire v_S_9458_out0;
wire v_S_9459_out0;
wire v_S_9460_out0;
wire v_S_9461_out0;
wire v_S_9462_out0;
wire v_S_9463_out0;
wire v_S_9464_out0;
wire v_S_9465_out0;
wire v_S_9466_out0;
wire v_S_9467_out0;
wire v_S_9468_out0;
wire v_S_9469_out0;
wire v_S_9470_out0;
wire v_S_9471_out0;
wire v_S_9472_out0;
wire v_S_9473_out0;
wire v_S_9474_out0;
wire v_S_9475_out0;
wire v_S_9476_out0;
wire v_S_9477_out0;
wire v_S_9478_out0;
wire v_S_9479_out0;
wire v_S_9480_out0;
wire v_S_9481_out0;
wire v_S_9482_out0;
wire v_S_9483_out0;
wire v_S_9484_out0;
wire v_S_9485_out0;
wire v_S_9486_out0;
wire v_S_9487_out0;
wire v_S_9488_out0;
wire v_S_9489_out0;
wire v_S_9490_out0;
wire v_S_9491_out0;
wire v_S_9492_out0;
wire v_S_9493_out0;
wire v_S_9494_out0;
wire v_S_9495_out0;
wire v_S_9496_out0;
wire v_S_9497_out0;
wire v_S_9498_out0;
wire v_S_9499_out0;
wire v_S_9500_out0;
wire v_S_9501_out0;
wire v_S_9502_out0;
wire v_S_9503_out0;
wire v_S_9504_out0;
wire v_S_9505_out0;
wire v_S_9506_out0;
wire v_S_9507_out0;
wire v_S_9508_out0;
wire v_S_9509_out0;
wire v_S_9510_out0;
wire v_S_9511_out0;
wire v_S_9512_out0;
wire v_S_9513_out0;
wire v_S_9514_out0;
wire v_S_9515_out0;
wire v_S_9516_out0;
wire v_S_9517_out0;
wire v_S_9518_out0;
wire v_S_9519_out0;
wire v_S_9520_out0;
wire v_S_9521_out0;
wire v_S_9522_out0;
wire v_S_9523_out0;
wire v_S_9524_out0;
wire v_S_9525_out0;
wire v_S_9526_out0;
wire v_S_9527_out0;
wire v_S_9528_out0;
wire v_S_9529_out0;
wire v_S_9530_out0;
wire v_S_9531_out0;
wire v_S_9532_out0;
wire v_S_9533_out0;
wire v_S_9534_out0;
wire v_S_9535_out0;
wire v_S_9536_out0;
wire v_S_9537_out0;
wire v_S_9538_out0;
wire v_S_9539_out0;
wire v_S_9540_out0;
wire v_S_9541_out0;
wire v_S_9542_out0;
wire v_S_9543_out0;
wire v_S_9544_out0;
wire v_S_9545_out0;
wire v_S_9546_out0;
wire v_S_9547_out0;
wire v_S_9548_out0;
wire v_S_9549_out0;
wire v_S_9550_out0;
wire v_S_9551_out0;
wire v_S_9552_out0;
wire v_S_9553_out0;
wire v_S_9554_out0;
wire v_S_9555_out0;
wire v_S_9556_out0;
wire v_S_9557_out0;
wire v_S_9558_out0;
wire v_S_9559_out0;
wire v_S_9560_out0;
wire v_S_9561_out0;
wire v_S_9562_out0;
wire v_S_9563_out0;
wire v_S_9564_out0;
wire v_S_9565_out0;
wire v_S_9566_out0;
wire v_S_9567_out0;
wire v_S_9568_out0;
wire v_S_9569_out0;
wire v_S_9570_out0;
wire v_S_9571_out0;
wire v_S_9572_out0;
wire v_S_9573_out0;
wire v_S_9574_out0;
wire v_S_9575_out0;
wire v_S_9576_out0;
wire v_S_9577_out0;
wire v_S_9578_out0;
wire v_S_9579_out0;
wire v_S_9580_out0;
wire v_S_9581_out0;
wire v_S_9582_out0;
wire v_S_9583_out0;
wire v_S_9584_out0;
wire v_S_9585_out0;
wire v_S_9586_out0;
wire v_S_9587_out0;
wire v_S_9588_out0;
wire v_S_9589_out0;
wire v_S_9590_out0;
wire v_S_9591_out0;
wire v_S_9592_out0;
wire v_S_9593_out0;
wire v_S_9594_out0;
wire v_S_9595_out0;
wire v_S_9596_out0;
wire v_S_9597_out0;
wire v_S_9598_out0;
wire v_S_9599_out0;
wire v_S_9600_out0;
wire v_S_9601_out0;
wire v_S_9602_out0;
wire v_S_9603_out0;
wire v_S_9604_out0;
wire v_S_9605_out0;
wire v_S_9606_out0;
wire v_S_9607_out0;
wire v_S_9608_out0;
wire v_S_9609_out0;
wire v_S_9610_out0;
wire v_S_9611_out0;
wire v_S_9612_out0;
wire v_S_9613_out0;
wire v_S_9614_out0;
wire v_S_9615_out0;
wire v_S_9616_out0;
wire v_S_9617_out0;
wire v_S_9618_out0;
wire v_S_9619_out0;
wire v_S_9620_out0;
wire v_S_9621_out0;
wire v_S_9622_out0;
wire v_S_9623_out0;
wire v_S_9624_out0;
wire v_S_9625_out0;
wire v_S_9626_out0;
wire v_S_9627_out0;
wire v_S_9628_out0;
wire v_S_9629_out0;
wire v_S_9630_out0;
wire v_S_9631_out0;
wire v_S_9632_out0;
wire v_S_9633_out0;
wire v_S_9634_out0;
wire v_S_9635_out0;
wire v_S_9636_out0;
wire v_S_9637_out0;
wire v_S_9638_out0;
wire v_S_9639_out0;
wire v_S_9640_out0;
wire v_S_9641_out0;
wire v_S_9642_out0;
wire v_S_9643_out0;
wire v_S_9644_out0;
wire v_S_9645_out0;
wire v_S_9646_out0;
wire v_S_9647_out0;
wire v_S_9648_out0;
wire v_S_9649_out0;
wire v_S_9650_out0;
wire v_S_9651_out0;
wire v_S_9652_out0;
wire v_S_9653_out0;
wire v_S_9654_out0;
wire v_S_9655_out0;
wire v_S_9656_out0;
wire v_S_9657_out0;
wire v_S_9658_out0;
wire v_S_9659_out0;
wire v_S_9660_out0;
wire v_S_9661_out0;
wire v_S_9662_out0;
wire v_S_9663_out0;
wire v_S_9664_out0;
wire v_S_9665_out0;
wire v_S_9666_out0;
wire v_S_9667_out0;
wire v_S_9668_out0;
wire v_S_9669_out0;
wire v_S_9670_out0;
wire v_S_9671_out0;
wire v_S_9672_out0;
wire v_S_9673_out0;
wire v_S_9674_out0;
wire v_S_9675_out0;
wire v_S_9676_out0;
wire v_S_9677_out0;
wire v_S_9678_out0;
wire v_S_9679_out0;
wire v_S_9680_out0;
wire v_S_9681_out0;
wire v_S_9682_out0;
wire v_S_9683_out0;
wire v_S_9684_out0;
wire v_S_9685_out0;
wire v_S_9686_out0;
wire v_S_9687_out0;
wire v_S_9688_out0;
wire v_S_9689_out0;
wire v_S_9690_out0;
wire v_S_9691_out0;
wire v_S_9692_out0;
wire v_S_9693_out0;
wire v_S_9694_out0;
wire v_S_9695_out0;
wire v_S_9696_out0;
wire v_S_9697_out0;
wire v_S_9698_out0;
wire v_S_9699_out0;
wire v_S_9700_out0;
wire v_S_9701_out0;
wire v_S_9702_out0;
wire v_S_9703_out0;
wire v_S_9704_out0;
wire v_S_9705_out0;
wire v_S_9706_out0;
wire v_S_9707_out0;
wire v_S_9708_out0;
wire v_S_9709_out0;
wire v_S_9710_out0;
wire v_S_9711_out0;
wire v_S_9712_out0;
wire v_S_9713_out0;
wire v_S_9714_out0;
wire v_S_9715_out0;
wire v_S_9716_out0;
wire v_S_9717_out0;
wire v_S_9718_out0;
wire v_S_9719_out0;
wire v_S_9720_out0;
wire v_S_9721_out0;
wire v_S_9722_out0;
wire v_S_9723_out0;
wire v_S_9724_out0;
wire v_S_9725_out0;
wire v_S_9726_out0;
wire v_S_9727_out0;
wire v_S_9728_out0;
wire v_S_9729_out0;
wire v_S_9730_out0;
wire v_S_9731_out0;
wire v_S_9732_out0;
wire v_S_9733_out0;
wire v_S_9734_out0;
wire v_S_9735_out0;
wire v_S_9736_out0;
wire v_S_9737_out0;
wire v_S_9738_out0;
wire v_S_9739_out0;
wire v_S_9740_out0;
wire v_S_9741_out0;
wire v_S_9742_out0;
wire v_S_9743_out0;
wire v_S_9744_out0;
wire v_S_9745_out0;
wire v_S_9746_out0;
wire v_S_9747_out0;
wire v_S_9748_out0;
wire v_S_9749_out0;
wire v_S_9750_out0;
wire v_S_9751_out0;
wire v_S_9752_out0;
wire v_S_9753_out0;
wire v_S_9754_out0;
wire v_S_9755_out0;
wire v_S_9756_out0;
wire v_S_9757_out0;
wire v_S_9758_out0;
wire v_S_9759_out0;
wire v_S_9760_out0;
wire v_S_9761_out0;
wire v_S_9762_out0;
wire v_S_9763_out0;
wire v_S_9764_out0;
wire v_S_9765_out0;
wire v_S_9766_out0;
wire v_S_9767_out0;
wire v_S_9768_out0;
wire v_S_9769_out0;
wire v_S_9770_out0;
wire v_S_9771_out0;
wire v_S_9772_out0;
wire v_S_9773_out0;
wire v_S_9774_out0;
wire v_S_9775_out0;
wire v_S_9776_out0;
wire v_S_9777_out0;
wire v_S_9778_out0;
wire v_S_9779_out0;
wire v_S_9780_out0;
wire v_S_9781_out0;
wire v_S_9782_out0;
wire v_S_9783_out0;
wire v_S_9784_out0;
wire v_S_9785_out0;
wire v_S_9786_out0;
wire v_S_9787_out0;
wire v_S_9788_out0;
wire v_S_9789_out0;
wire v_S_9790_out0;
wire v_TRANSMIT_INSTRUCTION_1713_out0;
wire v_TST_3819_out0;
wire v_TST_3820_out0;
wire v_TST_409_out0;
wire v_TST_410_out0;
wire v_TST_8735_out0;
wire v_TST_8736_out0;
wire v_TX_INSTRUCTION0_1762_out0;
wire v_TX_INSTRUCTION1_1169_out0;
wire v_TX_INSTRUCTION_10501_out0;
wire v_TX_INSTRUCTION_13631_out0;
wire v_TX_INSTRUCTION_13659_out0;
wire v_TX_INSTRUCTION_13660_out0;
wire v_TX_INSTRUCTION_2825_out0;
wire v_TX_INSTRUCTION_453_out0;
wire v_TX_INSTRUCTION_62_out0;
wire v_TX_INSTRUCTION_63_out0;
wire v_TX_INSTRUCTION_6875_out0;
wire v_TX_INSTRUCTION_7012_out0;
wire v_TX_INSTRUCTION_7013_out0;
wire v_TX_INSTUCTION0_228_out0;
wire v_TX_INSTUCTION1_4859_out0;
wire v_TX_INST_10827_out0;
wire v_TX_INST_10828_out0;
wire v_TX_INST_11239_out0;
wire v_TX_IN_PROGRESS_13634_out0;
wire v_TX_IN_PROGRESS_235_out0;
wire v_TX_OVERFLOW_10481_out0;
wire v_TX_OVERFLOW_13294_out0;
wire v_TX_OVERFLOW_500_out0;
wire v_TX_PROGRESS_8645_out0;
wire v_TX_inst0_608_out0;
wire v_UART_10516_out0;
wire v_UART_10517_out0;
wire v_UART_10825_out0;
wire v_UART_10826_out0;
wire v_UART_11128_out0;
wire v_UART_11129_out0;
wire v_UART_1823_out0;
wire v_UART_1824_out0;
wire v_UART_3893_out0;
wire v_UART_3894_out0;
wire v_UNDERFLOW_6916_out0;
wire v_UNDERFLOW_6917_out0;
wire v_UNNOTUSED_11220_out0;
wire v_UNNOTUSED_11221_out0;
wire v_UNUSED1_3016_out0;
wire v_UNUSED1_3017_out0;
wire v_UNUSED1_3220_out0;
wire v_UNUSED2_2193_out0;
wire v_UNUSED2_2194_out0;
wire v_UNUSED2_2424_out0;
wire v_UNUSED3_1681_out0;
wire v_UNUSED_123_out0;
wire v_UNUSED_339_out0;
wire v_UNUSED_340_out0;
wire v_U_10469_out0;
wire v_U_10470_out0;
wire v_WEN0_13300_out0;
wire v_WEN0_2588_out0;
wire v_WEN0_2646_out0;
wire v_WEN1_7716_out0;
wire v_WEN1_8763_out0;
wire v_WEN3_1690_out0;
wire v_WEN3_1691_out0;
wire v_WENALU_10866_out0;
wire v_WENALU_10867_out0;
wire v_WENALU_8659_out0;
wire v_WENALU_8660_out0;
wire v_WENLDST_13755_out0;
wire v_WENLDST_13756_out0;
wire v_WENLDST_2682_out0;
wire v_WENLDST_2683_out0;
wire v_WENLS_11260_out0;
wire v_WENLS_11261_out0;
wire v_WENLS_600_out0;
wire v_WENLS_601_out0;
wire v_WENMULTI_11206_out0;
wire v_WENMULTI_11207_out0;
wire v_WENRAM_2326_out0;
wire v_WENRAM_2327_out0;
wire v_WENRAM_4650_out0;
wire v_WENRAM_4651_out0;
wire v_WEN_11038_out0;
wire v_WEN_11039_out0;
wire v_WEN_2154_out0;
wire v_WEN_2765_out0;
wire v_WEN_2766_out0;
wire v_WEN_3204_out0;
wire v_WEN_MULTI_10381_out0;
wire v_WEN_MULTI_10382_out0;
wire v_WEN_MULTI_2388_out0;
wire v_WEN_MULTI_2389_out0;
wire v_WEN_MULTI_35_out0;
wire v_WEN_MULTI_36_out0;
wire v_WEN_RAM_7079_out0;
wire v_WEN_RAM_7080_out0;
wire v_WRITE_EN_13653_out0;
wire v_WRITE_EN_13654_out0;
wire v_WWNELS0_385_out0;
wire v_WWNELS1_47_out0;
wire v_W_EN_6878_out0;
wire v_W_EN_6879_out0;
wire v_Wen1_10312_out0;
wire v__0_out0;
wire v__10377_out0;
wire v__10378_out0;
wire v__10379_out0;
wire v__10380_out0;
wire v__10385_out0;
wire v__10386_out0;
wire v__10387_out0;
wire v__10388_out0;
wire v__10409_out0;
wire v__10410_out0;
wire v__10411_out0;
wire v__10412_out0;
wire v__10413_out0;
wire v__10414_out0;
wire v__10415_out0;
wire v__10416_out0;
wire v__10417_out0;
wire v__10418_out0;
wire v__10419_out0;
wire v__10420_out0;
wire v__10421_out0;
wire v__10422_out0;
wire v__10423_out0;
wire v__10424_out0;
wire v__10425_out0;
wire v__10426_out0;
wire v__10427_out0;
wire v__10428_out0;
wire v__10429_out0;
wire v__10430_out0;
wire v__10431_out0;
wire v__10432_out0;
wire v__10433_out0;
wire v__10434_out0;
wire v__10435_out0;
wire v__10436_out0;
wire v__10437_out0;
wire v__10438_out0;
wire v__10472_out0;
wire v__10473_out0;
wire v__10479_out0;
wire v__10480_out0;
wire v__10490_out1;
wire v__10491_out1;
wire v__10536_out0;
wire v__10537_out0;
wire v__10538_out0;
wire v__10539_out0;
wire v__10695_out0;
wire v__10696_out0;
wire v__10697_out0;
wire v__10698_out0;
wire v__10717_out0;
wire v__10718_out0;
wire v__10719_out0;
wire v__10720_out0;
wire v__10721_out0;
wire v__10722_out0;
wire v__10723_out0;
wire v__10724_out0;
wire v__10725_out0;
wire v__10726_out0;
wire v__10727_out0;
wire v__10728_out0;
wire v__10729_out0;
wire v__10730_out0;
wire v__10731_out0;
wire v__10732_out0;
wire v__10733_out0;
wire v__10734_out0;
wire v__10735_out0;
wire v__10736_out0;
wire v__10737_out0;
wire v__10738_out0;
wire v__10739_out0;
wire v__10740_out0;
wire v__10741_out0;
wire v__10742_out0;
wire v__10743_out0;
wire v__10744_out0;
wire v__10745_out0;
wire v__10746_out0;
wire v__10747_out0;
wire v__10748_out0;
wire v__10777_out0;
wire v__10778_out0;
wire v__10779_out0;
wire v__10780_out0;
wire v__10785_out0;
wire v__10786_out0;
wire v__10808_out0;
wire v__10809_out0;
wire v__10823_out0;
wire v__10824_out0;
wire v__10862_out0;
wire v__10863_out0;
wire v__10864_out0;
wire v__10865_out0;
wire v__10868_out1;
wire v__10869_out1;
wire v__10874_out0;
wire v__10875_out0;
wire v__10876_out0;
wire v__10877_out0;
wire v__10878_out0;
wire v__10879_out0;
wire v__10880_out0;
wire v__10881_out0;
wire v__10882_out0;
wire v__10883_out0;
wire v__10884_out0;
wire v__10885_out0;
wire v__10886_out0;
wire v__10887_out0;
wire v__10888_out0;
wire v__10889_out0;
wire v__10890_out0;
wire v__10891_out0;
wire v__10892_out0;
wire v__10893_out0;
wire v__10894_out0;
wire v__10895_out0;
wire v__10896_out0;
wire v__10897_out0;
wire v__10898_out0;
wire v__10899_out0;
wire v__10900_out0;
wire v__10901_out0;
wire v__10902_out0;
wire v__10903_out0;
wire v__10910_out0;
wire v__10911_out0;
wire v__11001_out0;
wire v__11002_out0;
wire v__11003_out0;
wire v__11004_out0;
wire v__11005_out0;
wire v__11006_out0;
wire v__11007_out0;
wire v__11008_out0;
wire v__11009_out0;
wire v__11010_out0;
wire v__11011_out0;
wire v__11012_out0;
wire v__11013_out0;
wire v__11014_out0;
wire v__11015_out0;
wire v__11016_out0;
wire v__11017_out0;
wire v__11018_out0;
wire v__11019_out0;
wire v__11020_out0;
wire v__11021_out0;
wire v__11022_out0;
wire v__11023_out0;
wire v__11024_out0;
wire v__11025_out0;
wire v__11026_out0;
wire v__11027_out0;
wire v__11028_out0;
wire v__11029_out0;
wire v__11030_out0;
wire v__11098_out0;
wire v__11099_out0;
wire v__11100_out0;
wire v__11101_out0;
wire v__11102_out0;
wire v__11103_out0;
wire v__11104_out0;
wire v__11105_out0;
wire v__11106_out0;
wire v__11107_out0;
wire v__11108_out0;
wire v__11109_out0;
wire v__11110_out0;
wire v__11111_out0;
wire v__11112_out0;
wire v__11113_out0;
wire v__11114_out0;
wire v__11115_out0;
wire v__11116_out0;
wire v__11117_out0;
wire v__11118_out0;
wire v__11119_out0;
wire v__11120_out0;
wire v__11121_out0;
wire v__11122_out0;
wire v__11123_out0;
wire v__11124_out0;
wire v__11125_out0;
wire v__11126_out0;
wire v__11127_out0;
wire v__11149_out0;
wire v__11150_out0;
wire v__11151_out0;
wire v__11152_out0;
wire v__11212_out0;
wire v__11213_out0;
wire v__11242_out0;
wire v__11243_out0;
wire v__11294_out1;
wire v__11295_out1;
wire v__1176_out0;
wire v__1177_out0;
wire v__1193_out0;
wire v__1194_out0;
wire v__13251_out0;
wire v__13252_out0;
wire v__13384_out0;
wire v__13385_out0;
wire v__13386_out0;
wire v__13387_out0;
wire v__13392_out0;
wire v__13393_out0;
wire v__13396_out0;
wire v__13397_out0;
wire v__13399_out0;
wire v__13400_out0;
wire v__13401_out0;
wire v__13402_out0;
wire v__13403_out0;
wire v__13404_out0;
wire v__13405_out0;
wire v__13406_out0;
wire v__13407_out0;
wire v__13408_out0;
wire v__13409_out0;
wire v__13410_out0;
wire v__13411_out0;
wire v__13412_out0;
wire v__13413_out0;
wire v__13414_out0;
wire v__13415_out0;
wire v__13416_out0;
wire v__13417_out0;
wire v__13418_out0;
wire v__13419_out0;
wire v__13420_out0;
wire v__13421_out0;
wire v__13422_out0;
wire v__13423_out0;
wire v__13424_out0;
wire v__13425_out0;
wire v__13426_out0;
wire v__13427_out0;
wire v__13428_out0;
wire v__13435_out0;
wire v__13436_out0;
wire v__13448_out0;
wire v__13449_out0;
wire v__13450_out0;
wire v__13451_out0;
wire v__13452_out0;
wire v__13453_out0;
wire v__13454_out0;
wire v__13455_out0;
wire v__13456_out0;
wire v__13457_out0;
wire v__13458_out0;
wire v__13459_out0;
wire v__13460_out0;
wire v__13461_out0;
wire v__13462_out0;
wire v__13463_out0;
wire v__13464_out0;
wire v__13465_out0;
wire v__13466_out0;
wire v__13467_out0;
wire v__13468_out0;
wire v__13469_out0;
wire v__13470_out0;
wire v__13471_out0;
wire v__13472_out0;
wire v__13473_out0;
wire v__13474_out0;
wire v__13475_out0;
wire v__13476_out0;
wire v__13477_out0;
wire v__13512_out0;
wire v__13513_out0;
wire v__13514_out0;
wire v__13515_out0;
wire v__13552_out0;
wire v__13553_out0;
wire v__13554_out0;
wire v__13555_out0;
wire v__13562_out0;
wire v__13563_out0;
wire v__13601_out0;
wire v__13602_out0;
wire v__13627_out0;
wire v__13628_out0;
wire v__13629_out0;
wire v__13630_out0;
wire v__13715_out0;
wire v__13716_out0;
wire v__13717_out0;
wire v__13718_out0;
wire v__13719_out0;
wire v__13720_out0;
wire v__13721_out0;
wire v__13722_out0;
wire v__13723_out0;
wire v__13724_out0;
wire v__13725_out0;
wire v__13726_out0;
wire v__13727_out0;
wire v__13728_out0;
wire v__13729_out0;
wire v__13730_out0;
wire v__13731_out0;
wire v__13732_out0;
wire v__13733_out0;
wire v__13734_out0;
wire v__13735_out0;
wire v__13736_out0;
wire v__13737_out0;
wire v__13738_out0;
wire v__13739_out0;
wire v__13740_out0;
wire v__13741_out0;
wire v__13742_out0;
wire v__13743_out0;
wire v__13744_out0;
wire v__1692_out0;
wire v__1693_out0;
wire v__1694_out0;
wire v__1695_out0;
wire v__171_out0;
wire v__1722_out0;
wire v__1723_out0;
wire v__1724_out0;
wire v__1725_out0;
wire v__1728_out0;
wire v__1729_out0;
wire v__172_out0;
wire v__1747_out0;
wire v__1748_out0;
wire v__1749_out0;
wire v__1750_out0;
wire v__1773_out0;
wire v__1774_out0;
wire v__1775_out0;
wire v__1776_out0;
wire v__1777_out0;
wire v__1778_out0;
wire v__1779_out0;
wire v__1780_out0;
wire v__1781_out0;
wire v__1782_out0;
wire v__1783_out0;
wire v__1784_out0;
wire v__1785_out0;
wire v__1786_out0;
wire v__1787_out0;
wire v__1788_out0;
wire v__1789_out0;
wire v__1790_out0;
wire v__1791_out0;
wire v__1792_out0;
wire v__1793_out0;
wire v__1794_out0;
wire v__1795_out0;
wire v__1796_out0;
wire v__1797_out0;
wire v__1798_out0;
wire v__1799_out0;
wire v__179_out0;
wire v__1800_out0;
wire v__1801_out0;
wire v__1802_out0;
wire v__180_out0;
wire v__186_out0;
wire v__1875_out0;
wire v__1876_out0;
wire v__187_out0;
wire v__1893_out0;
wire v__1894_out0;
wire v__1895_out0;
wire v__1896_out0;
wire v__1904_out0;
wire v__1905_out0;
wire v__192_out0;
wire v__193_out0;
wire v__194_out0;
wire v__195_out0;
wire v__1975_out0;
wire v__1976_out0;
wire v__1977_out0;
wire v__1978_out0;
wire v__1979_out0;
wire v__1980_out0;
wire v__1981_out0;
wire v__1982_out0;
wire v__1983_out0;
wire v__1984_out0;
wire v__1985_out0;
wire v__1986_out0;
wire v__1987_out0;
wire v__1988_out0;
wire v__1989_out0;
wire v__198_out0;
wire v__1990_out0;
wire v__1991_out0;
wire v__1992_out0;
wire v__1993_out0;
wire v__1994_out0;
wire v__1995_out0;
wire v__1996_out0;
wire v__1997_out0;
wire v__1998_out0;
wire v__1999_out0;
wire v__199_out0;
wire v__1_out0;
wire v__2000_out0;
wire v__2001_out0;
wire v__2002_out0;
wire v__2003_out0;
wire v__2004_out0;
wire v__2022_out0;
wire v__2023_out0;
wire v__2063_out0;
wire v__2064_out0;
wire v__2065_out0;
wire v__2066_out0;
wire v__2067_out0;
wire v__2068_out0;
wire v__2069_out0;
wire v__2070_out0;
wire v__2071_out0;
wire v__2072_out0;
wire v__2073_out0;
wire v__2074_out0;
wire v__2075_out0;
wire v__2076_out0;
wire v__2077_out0;
wire v__2078_out0;
wire v__2079_out0;
wire v__2080_out0;
wire v__2081_out0;
wire v__2082_out0;
wire v__2083_out0;
wire v__2084_out0;
wire v__2085_out0;
wire v__2086_out0;
wire v__2087_out0;
wire v__2088_out0;
wire v__2089_out0;
wire v__2090_out0;
wire v__2091_out0;
wire v__2092_out0;
wire v__2093_out0;
wire v__2094_out0;
wire v__2095_out0;
wire v__2096_out0;
wire v__2150_out0;
wire v__2151_out0;
wire v__2152_out0;
wire v__2153_out0;
wire v__2155_out0;
wire v__2156_out0;
wire v__2157_out0;
wire v__2158_out0;
wire v__2159_out0;
wire v__2160_out0;
wire v__2161_out0;
wire v__2162_out0;
wire v__2163_out0;
wire v__2164_out0;
wire v__2165_out0;
wire v__2166_out0;
wire v__2167_out0;
wire v__2168_out0;
wire v__2169_out0;
wire v__2170_out0;
wire v__2171_out0;
wire v__2172_out0;
wire v__2173_out0;
wire v__2174_out0;
wire v__2175_out0;
wire v__2176_out0;
wire v__2177_out0;
wire v__2178_out0;
wire v__2179_out0;
wire v__2180_out0;
wire v__2181_out0;
wire v__2182_out0;
wire v__2183_out0;
wire v__2184_out0;
wire v__2195_out0;
wire v__2196_out0;
wire v__2197_out0;
wire v__2198_out0;
wire v__2199_out0;
wire v__2200_out0;
wire v__2201_out0;
wire v__2202_out0;
wire v__2203_out0;
wire v__2204_out0;
wire v__2205_out0;
wire v__2206_out0;
wire v__2207_out0;
wire v__2208_out0;
wire v__2209_out0;
wire v__2210_out0;
wire v__2211_out0;
wire v__2212_out0;
wire v__2213_out0;
wire v__2214_out0;
wire v__2215_out0;
wire v__2216_out0;
wire v__2217_out0;
wire v__2218_out0;
wire v__2219_out0;
wire v__2220_out0;
wire v__2221_out0;
wire v__2222_out0;
wire v__2268_out0;
wire v__2269_out0;
wire v__2273_out0;
wire v__2274_out0;
wire v__2275_out0;
wire v__2276_out0;
wire v__2277_out0;
wire v__2278_out0;
wire v__2279_out0;
wire v__2280_out0;
wire v__2281_out0;
wire v__2282_out0;
wire v__2283_out0;
wire v__2284_out0;
wire v__2285_out0;
wire v__2286_out0;
wire v__2287_out0;
wire v__2288_out0;
wire v__2289_out0;
wire v__2290_out0;
wire v__2291_out0;
wire v__2292_out0;
wire v__2293_out0;
wire v__2294_out0;
wire v__2295_out0;
wire v__2296_out0;
wire v__2297_out0;
wire v__2298_out0;
wire v__2299_out0;
wire v__2300_out0;
wire v__2301_out0;
wire v__2302_out0;
wire v__2418_out0;
wire v__2419_out0;
wire v__2420_out0;
wire v__2421_out0;
wire v__2422_out0;
wire v__2423_out0;
wire v__2430_out0;
wire v__2431_out0;
wire v__2462_out0;
wire v__2463_out0;
wire v__2467_out0;
wire v__2468_out0;
wire v__2470_out0;
wire v__2471_out0;
wire v__2502_out0;
wire v__2503_out0;
wire v__2504_out0;
wire v__2505_out0;
wire v__2506_out0;
wire v__2507_out0;
wire v__2508_out0;
wire v__2509_out0;
wire v__2510_out0;
wire v__2511_out0;
wire v__2512_out0;
wire v__2513_out0;
wire v__2514_out0;
wire v__2515_out0;
wire v__2516_out0;
wire v__2517_out0;
wire v__2518_out0;
wire v__2519_out0;
wire v__2520_out0;
wire v__2521_out0;
wire v__2522_out0;
wire v__2523_out0;
wire v__2524_out0;
wire v__2525_out0;
wire v__2526_out0;
wire v__2527_out0;
wire v__2528_out0;
wire v__2529_out0;
wire v__2530_out0;
wire v__2531_out0;
wire v__2692_out0;
wire v__2693_out0;
wire v__2726_out0;
wire v__2727_out0;
wire v__2728_out0;
wire v__2729_out0;
wire v__2730_out0;
wire v__2731_out0;
wire v__2732_out0;
wire v__2733_out0;
wire v__2734_out0;
wire v__2735_out0;
wire v__2736_out0;
wire v__2737_out0;
wire v__2738_out0;
wire v__2739_out0;
wire v__2740_out0;
wire v__2741_out0;
wire v__2742_out0;
wire v__2743_out0;
wire v__2744_out0;
wire v__2745_out0;
wire v__2746_out0;
wire v__2747_out0;
wire v__2748_out0;
wire v__2749_out0;
wire v__2750_out0;
wire v__2751_out0;
wire v__2752_out0;
wire v__2753_out0;
wire v__2754_out0;
wire v__2755_out0;
wire v__2760_out0;
wire v__2761_out0;
wire v__2762_out0;
wire v__2763_out0;
wire v__2831_out0;
wire v__2831_out1;
wire v__2832_out0;
wire v__2832_out1;
wire v__2860_out0;
wire v__2861_out0;
wire v__2875_out0;
wire v__2876_out0;
wire v__2877_out0;
wire v__2878_out0;
wire v__2879_out0;
wire v__287_out0;
wire v__2880_out0;
wire v__2881_out0;
wire v__2882_out0;
wire v__2889_out0;
wire v__288_out0;
wire v__2890_out0;
wire v__2943_out0;
wire v__2944_out0;
wire v__2959_out0;
wire v__2973_out0;
wire v__2974_out0;
wire v__2983_out0;
wire v__2983_out1;
wire v__2984_out0;
wire v__2985_out0;
wire v__2986_out0;
wire v__2987_out0;
wire v__2988_out0;
wire v__2989_out0;
wire v__2990_out0;
wire v__2991_out0;
wire v__2992_out0;
wire v__2993_out0;
wire v__2994_out0;
wire v__2995_out0;
wire v__2996_out0;
wire v__2997_out0;
wire v__2998_out0;
wire v__2999_out0;
wire v__2_out0;
wire v__3000_out0;
wire v__3001_out0;
wire v__3002_out0;
wire v__3003_out0;
wire v__3004_out0;
wire v__3005_out0;
wire v__3006_out0;
wire v__3007_out0;
wire v__3008_out0;
wire v__3009_out0;
wire v__3010_out0;
wire v__3011_out0;
wire v__3012_out0;
wire v__3013_out0;
wire v__3014_out0;
wire v__3015_out0;
wire v__3051_out0;
wire v__3052_out0;
wire v__3053_out0;
wire v__3054_out0;
wire v__3055_out0;
wire v__3056_out0;
wire v__3057_out0;
wire v__3058_out0;
wire v__3059_out0;
wire v__3060_out0;
wire v__3061_out0;
wire v__3062_out0;
wire v__3063_out0;
wire v__3064_out0;
wire v__3065_out0;
wire v__3066_out0;
wire v__3067_out0;
wire v__3068_out0;
wire v__3069_out0;
wire v__3070_out0;
wire v__3071_out0;
wire v__3072_out0;
wire v__3073_out0;
wire v__3074_out0;
wire v__3075_out0;
wire v__3076_out0;
wire v__3077_out0;
wire v__3078_out0;
wire v__3079_out0;
wire v__3080_out0;
wire v__3085_out0;
wire v__3086_out0;
wire v__3087_out0;
wire v__3088_out0;
wire v__3089_out0;
wire v__3090_out0;
wire v__3091_out0;
wire v__3092_out0;
wire v__3093_out0;
wire v__3094_out0;
wire v__3095_out0;
wire v__3096_out0;
wire v__3097_out0;
wire v__3098_out0;
wire v__3099_out0;
wire v__3100_out0;
wire v__3101_out0;
wire v__3102_out0;
wire v__3103_out0;
wire v__3104_out0;
wire v__3105_out0;
wire v__3106_out0;
wire v__3107_out0;
wire v__3108_out0;
wire v__3109_out0;
wire v__3110_out0;
wire v__3111_out0;
wire v__3112_out0;
wire v__3113_out0;
wire v__3114_out0;
wire v__3119_out0;
wire v__3120_out0;
wire v__3121_out0;
wire v__3122_out0;
wire v__3123_out0;
wire v__3124_out0;
wire v__3139_out0;
wire v__3140_out0;
wire v__3141_out0;
wire v__3142_out0;
wire v__3143_out0;
wire v__3144_out0;
wire v__3145_out0;
wire v__3146_out0;
wire v__3147_out0;
wire v__3148_out0;
wire v__3149_out0;
wire v__3150_out0;
wire v__3151_out0;
wire v__3152_out0;
wire v__3153_out0;
wire v__3154_out0;
wire v__3155_out0;
wire v__3156_out0;
wire v__3157_out0;
wire v__3158_out0;
wire v__3159_out0;
wire v__3160_out0;
wire v__3161_out0;
wire v__3162_out0;
wire v__3163_out0;
wire v__3164_out0;
wire v__3165_out0;
wire v__3166_out0;
wire v__3167_out0;
wire v__3168_out0;
wire v__3180_out0;
wire v__3181_out0;
wire v__3199_out0;
wire v__3200_out0;
wire v__321_out0;
wire v__322_out0;
wire v__3237_out0;
wire v__3238_out0;
wire v__323_out0;
wire v__3247_out0;
wire v__3248_out0;
wire v__3249_out0;
wire v__324_out0;
wire v__3250_out0;
wire v__3266_out0;
wire v__3267_out0;
wire v__3270_out0;
wire v__3271_out0;
wire v__3282_out0;
wire v__3283_out0;
wire v__3284_out0;
wire v__3285_out0;
wire v__329_out0;
wire v__330_out0;
wire v__331_out0;
wire v__332_out0;
wire v__37_out0;
wire v__3803_out0;
wire v__3804_out0;
wire v__3823_out0;
wire v__3824_out0;
wire v__3825_out0;
wire v__3826_out0;
wire v__3827_out0;
wire v__3828_out0;
wire v__3829_out0;
wire v__3830_out0;
wire v__3831_out0;
wire v__3832_out0;
wire v__3833_out0;
wire v__3834_out0;
wire v__3835_out0;
wire v__3836_out0;
wire v__3837_out0;
wire v__3838_out0;
wire v__3839_out0;
wire v__3840_out0;
wire v__3841_out0;
wire v__3842_out0;
wire v__3843_out0;
wire v__3844_out0;
wire v__3845_out0;
wire v__3846_out0;
wire v__3847_out0;
wire v__3848_out0;
wire v__3849_out0;
wire v__3850_out0;
wire v__3851_out0;
wire v__3852_out0;
wire v__3861_out0;
wire v__3862_out0;
wire v__3863_out0;
wire v__3864_out0;
wire v__3865_out0;
wire v__3866_out0;
wire v__3867_out0;
wire v__3868_out0;
wire v__3869_out0;
wire v__3870_out0;
wire v__3871_out0;
wire v__3872_out0;
wire v__3873_out0;
wire v__3874_out0;
wire v__3875_out0;
wire v__3876_out0;
wire v__3877_out0;
wire v__3878_out0;
wire v__3879_out0;
wire v__3880_out0;
wire v__3881_out0;
wire v__3882_out0;
wire v__3883_out0;
wire v__3884_out0;
wire v__3885_out0;
wire v__3886_out0;
wire v__3887_out0;
wire v__3888_out0;
wire v__3889_out0;
wire v__3890_out0;
wire v__38_out0;
wire v__3907_out0;
wire v__3908_out0;
wire v__3910_out0;
wire v__3911_out0;
wire v__3912_out0;
wire v__3913_out0;
wire v__3914_out0;
wire v__3915_out0;
wire v__3916_out0;
wire v__3917_out0;
wire v__3918_out0;
wire v__3919_out0;
wire v__3920_out0;
wire v__3921_out0;
wire v__3922_out0;
wire v__3923_out0;
wire v__3924_out0;
wire v__3925_out0;
wire v__3926_out0;
wire v__3927_out0;
wire v__3928_out0;
wire v__3929_out0;
wire v__3930_out0;
wire v__3931_out0;
wire v__3932_out0;
wire v__3933_out0;
wire v__3934_out0;
wire v__3935_out0;
wire v__3936_out0;
wire v__3937_out0;
wire v__3938_out0;
wire v__3939_out0;
wire v__3961_out0;
wire v__3962_out0;
wire v__3963_out0;
wire v__3964_out0;
wire v__3965_out0;
wire v__3966_out0;
wire v__3967_out0;
wire v__3968_out0;
wire v__3969_out0;
wire v__3970_out0;
wire v__3971_out0;
wire v__3972_out0;
wire v__3973_out0;
wire v__3974_out0;
wire v__3975_out0;
wire v__3976_out0;
wire v__3977_out0;
wire v__3978_out0;
wire v__3979_out0;
wire v__3980_out0;
wire v__3981_out0;
wire v__3982_out0;
wire v__3983_out0;
wire v__3984_out0;
wire v__3985_out0;
wire v__3986_out0;
wire v__3987_out0;
wire v__3988_out0;
wire v__3989_out0;
wire v__3990_out0;
wire v__3_out0;
wire v__413_out0;
wire v__414_out0;
wire v__437_out0;
wire v__438_out0;
wire v__4526_out1;
wire v__4527_out1;
wire v__4597_out0;
wire v__4598_out0;
wire v__4599_out0;
wire v__4600_out0;
wire v__4605_out0;
wire v__4605_out1;
wire v__4606_out0;
wire v__4606_out1;
wire v__4610_out0;
wire v__4611_out0;
wire v__468_out0;
wire v__469_out0;
wire v__470_out0;
wire v__4711_out0;
wire v__4712_out0;
wire v__4713_out0;
wire v__4714_out0;
wire v__471_out0;
wire v__472_out0;
wire v__473_out0;
wire v__474_out0;
wire v__475_out0;
wire v__476_out0;
wire v__477_out0;
wire v__478_out0;
wire v__479_out0;
wire v__480_out0;
wire v__4812_out0;
wire v__4813_out0;
wire v__4814_out0;
wire v__4815_out0;
wire v__481_out0;
wire v__482_out0;
wire v__4831_out1;
wire v__4832_out1;
wire v__4833_out0;
wire v__4834_out0;
wire v__4837_out0;
wire v__4838_out0;
wire v__483_out0;
wire v__484_out0;
wire v__4856_out0;
wire v__4857_out0;
wire v__485_out0;
wire v__486_out0;
wire v__487_out0;
wire v__488_out0;
wire v__489_out0;
wire v__490_out0;
wire v__491_out0;
wire v__492_out0;
wire v__493_out0;
wire v__494_out0;
wire v__495_out0;
wire v__496_out0;
wire v__497_out0;
wire v__503_out0;
wire v__504_out0;
wire v__505_out0;
wire v__506_out0;
wire v__507_out0;
wire v__508_out0;
wire v__509_out0;
wire v__510_out0;
wire v__511_out0;
wire v__512_out0;
wire v__513_out0;
wire v__514_out0;
wire v__515_out0;
wire v__516_out0;
wire v__517_out0;
wire v__518_out0;
wire v__519_out0;
wire v__520_out0;
wire v__521_out0;
wire v__522_out0;
wire v__523_out0;
wire v__524_out0;
wire v__525_out0;
wire v__526_out0;
wire v__527_out0;
wire v__528_out0;
wire v__529_out0;
wire v__530_out0;
wire v__531_out0;
wire v__532_out0;
wire v__568_out0;
wire v__569_out0;
wire v__570_out0;
wire v__571_out0;
wire v__572_out0;
wire v__573_out0;
wire v__574_out0;
wire v__575_out0;
wire v__576_out0;
wire v__577_out0;
wire v__578_out0;
wire v__579_out0;
wire v__580_out0;
wire v__581_out0;
wire v__582_out0;
wire v__5832_out0;
wire v__5832_out1;
wire v__5833_out0;
wire v__5833_out1;
wire v__583_out0;
wire v__584_out0;
wire v__585_out0;
wire v__5860_out0;
wire v__5860_out1;
wire v__586_out0;
wire v__587_out0;
wire v__588_out0;
wire v__589_out0;
wire v__590_out0;
wire v__591_out0;
wire v__592_out0;
wire v__593_out0;
wire v__594_out0;
wire v__595_out0;
wire v__596_out0;
wire v__597_out0;
wire v__60_out0;
wire v__61_out0;
wire v__6800_out0;
wire v__6801_out0;
wire v__6802_out0;
wire v__6803_out0;
wire v__6804_out0;
wire v__6805_out0;
wire v__6806_out0;
wire v__6807_out0;
wire v__6808_out0;
wire v__6809_out0;
wire v__6810_out0;
wire v__6811_out0;
wire v__6812_out0;
wire v__6813_out0;
wire v__6814_out0;
wire v__6815_out0;
wire v__6816_out0;
wire v__6817_out0;
wire v__6818_out0;
wire v__6819_out0;
wire v__6820_out0;
wire v__6821_out0;
wire v__6822_out0;
wire v__6823_out0;
wire v__6824_out0;
wire v__6825_out0;
wire v__6826_out0;
wire v__6827_out0;
wire v__6828_out0;
wire v__6829_out0;
wire v__6830_out0;
wire v__6831_out0;
wire v__6832_out0;
wire v__6833_out0;
wire v__6834_out0;
wire v__6835_out0;
wire v__6836_out0;
wire v__6837_out0;
wire v__6838_out0;
wire v__6839_out0;
wire v__6840_out0;
wire v__6841_out0;
wire v__6842_out0;
wire v__6843_out0;
wire v__6844_out0;
wire v__6845_out0;
wire v__6846_out0;
wire v__6847_out0;
wire v__6848_out0;
wire v__6849_out0;
wire v__6850_out0;
wire v__6851_out0;
wire v__6852_out0;
wire v__6853_out0;
wire v__6854_out0;
wire v__6855_out0;
wire v__6856_out0;
wire v__6857_out0;
wire v__6858_out0;
wire v__6859_out0;
wire v__6876_out0;
wire v__6876_out1;
wire v__6877_out0;
wire v__6877_out1;
wire v__7062_out1;
wire v__7063_out1;
wire v__7070_out0;
wire v__7071_out0;
wire v__7095_out0;
wire v__7096_out0;
wire v__7108_out0;
wire v__7109_out0;
wire v__7644_out0;
wire v__7645_out0;
wire v__7646_out0;
wire v__7647_out0;
wire v__7648_out0;
wire v__7649_out0;
wire v__7650_out0;
wire v__7651_out0;
wire v__7652_out0;
wire v__7653_out0;
wire v__7654_out0;
wire v__7655_out0;
wire v__7656_out0;
wire v__7657_out0;
wire v__7658_out0;
wire v__7659_out0;
wire v__7660_out0;
wire v__7661_out0;
wire v__7662_out0;
wire v__7663_out0;
wire v__7664_out0;
wire v__7665_out0;
wire v__7666_out0;
wire v__7667_out0;
wire v__7668_out0;
wire v__7669_out0;
wire v__7670_out0;
wire v__7671_out0;
wire v__7672_out0;
wire v__7673_out0;
wire v__77_out0;
wire v__78_out0;
wire v__79_out0;
wire v__80_out0;
wire v__8699_out0;
wire v__8700_out0;
wire v__8701_out0;
wire v__8702_out0;
wire v__8703_out0;
wire v__8704_out0;
wire v__8705_out0;
wire v__8706_out0;
wire v__8707_out0;
wire v__8708_out0;
wire v__8709_out0;
wire v__8710_out0;
wire v__8711_out0;
wire v__8712_out0;
wire v__8713_out0;
wire v__8714_out0;
wire v__8715_out0;
wire v__8716_out0;
wire v__8717_out0;
wire v__8718_out0;
wire v__8719_out0;
wire v__8720_out0;
wire v__8721_out0;
wire v__8722_out0;
wire v__8723_out0;
wire v__8724_out0;
wire v__8725_out0;
wire v__8726_out0;
wire v__8727_out0;
wire v__8728_out0;
wire v__8748_out0;
wire v__8749_out0;
wire v__8750_out0;
wire v__8751_out0;
wire v__8769_out0;
wire v__8770_out0;
wire v__8771_out0;
wire v__8772_out0;
wire v__8773_out0;
wire v__8774_out0;
wire v__8775_out0;
wire v__8776_out0;
wire v__8777_out0;
wire v__8778_out0;
wire v__8779_out0;
wire v__8780_out0;
wire v__8781_out0;
wire v__8782_out0;
wire v__8783_out0;
wire v__8784_out0;
wire v__8785_out0;
wire v__8786_out0;
wire v__8787_out0;
wire v__8788_out0;
wire v__8789_out0;
wire v__8790_out0;
wire v__8791_out0;
wire v__8792_out0;
wire v__8793_out0;
wire v__8794_out0;
wire v__8795_out0;
wire v__8796_out0;
wire v__8797_out0;
wire v__8798_out0;
wire v__8827_out0;
wire v__8828_out0;
wire v__8829_out0;
wire v__8830_out0;
wire v__8831_out0;
wire v__8832_out0;
wire v__8848_out0;
wire v__8849_out0;
wire v__8850_out0;
wire v__8851_out0;
wire v_byte_comp_10_2318_out0;
wire v_byte_comp_11_2645_out0;
wire v_byte_comp_1_6872_out0;
wire v_byte_comp_1_6923_out0;
wire v_byte_ready_5842_out0;
wire v_byte_ready_5843_out0;
wire v_done_receiving_10604_out0;
wire v_exec1ls_3341_out0;
wire v_exec1ls_3342_out0;
wire v_transmit_INSTRUCTION_2674_out0;
wire v_wen_ram_4595_out0;
wire v_wen_ram_4596_out0;

always @(posedge clk) v_FF1_48_out0 <= v_BYTE_READY_2852_out0;
always @(posedge clk) v_FF1_49_out0 <= v_BYTE_READY_2853_out0;
always @(posedge clk) v_FF6_112_out0 <= v_ENABLE_2651_out0 ? v_MUX5_13348_out0 : v_FF6_112_out0;
always @(posedge clk) v_REG1_432_out0 <= v_G19_10327_out0 ? v_MUX4_2658_out0 : v_REG1_432_out0;
always @(posedge clk) v_REG1_433_out0 <= v_G19_10328_out0 ? v_MUX4_2659_out0 : v_REG1_433_out0;
v_ROM1_462 I1 (v_ROM1_462_out0, v_REG1_7134_out0, clk);
always @(posedge clk) v_FF4_463_out0 <= v_ENABLE_2651_out0 ? v_MUX3_7140_out0 : v_FF4_463_out0;
v_RAM0_1680 I1 (v_RAM0_1680_out0, v_ADRESS_ins0_11169_out0, v_DATA_RAM_IN0_284_out0, v_DONE_RECEIVING_5857_out0, clk);
v_data_ram_1818 I1 (v_data_ram_1818_out0, v_ADRESS_8683_out0, v_DATA_2469_out0, v_WEN_2154_out0, clk);
always @(posedge clk) v_FF1_1955_out0 <= v_ENABLE_2651_out0 ? v_SEL1_13445_out0 : v_FF1_1955_out0;
always @(posedge clk) v_IHOLD_REGISTER_2013_out0 <= v_NORMAL_181_out0 ? v_RAM_OUT_1751_out0 : v_IHOLD_REGISTER_2013_out0;
always @(posedge clk) v_IHOLD_REGISTER_2014_out0 <= v_NORMAL_182_out0 ? v_RAM_OUT_1752_out0 : v_IHOLD_REGISTER_2014_out0;
always @(posedge clk) v_FF3_2016_out0 <= v_EN_7093_out0 ? v__4605_out0 : v_FF3_2016_out0;
always @(posedge clk) v_FF3_2017_out0 <= v_EN_7094_out0 ? v__4606_out0 : v_FF3_2017_out0;
always @(posedge clk) v_FF4_2106_out0 <= v_EN_7093_out0 ? v__4605_out1 : v_FF4_2106_out0;
always @(posedge clk) v_FF4_2107_out0 <= v_EN_7094_out0 ? v__4606_out1 : v_FF4_2107_out0;
always @(posedge clk) v_REG1_2314_out0 <= v_D1_8842_out1 ? v_DIN3_10310_out0 : v_REG1_2314_out0;
always @(posedge clk) v_REG1_2315_out0 <= v_D1_8843_out1 ? v_DIN3_10311_out0 : v_REG1_2315_out0;
always @(posedge clk) v_FF7_2670_out0 <= v_G24_10560_out0;
always @(posedge clk) v_FF7_2671_out0 <= v_G24_10561_out0;
always @(posedge clk) v_FF7_2672_out0 <= v_G24_10562_out0;
always @(posedge clk) v_FF7_2673_out0 <= v_G24_10563_out0;
always @(posedge clk) v_REG1_2677_out0 <= v_ENABLE_1757_out0 ? v__3040_out0 : v_REG1_2677_out0;
always @(posedge clk) v_FF2_2833_out0 <= v_ENABLE_2651_out0 ? v_MUX1_2625_out0 : v_FF2_2833_out0;
always @(posedge clk) v_FF1_4717_out0 <= v_EN_2919_out0 ? v_G1_2700_out0 : v_FF1_4717_out0;
always @(posedge clk) v_FF1_4718_out0 <= v_EN_2920_out0 ? v_G1_2701_out0 : v_FF1_4718_out0;
always @(posedge clk) v_FF1_4719_out0 <= v_EN_2921_out0 ? v_G1_2702_out0 : v_FF1_4719_out0;
always @(posedge clk) v_FF1_4720_out0 <= v_EN_2922_out0 ? v_G1_2703_out0 : v_FF1_4720_out0;
always @(posedge clk) v_FF1_4721_out0 <= v_EN_2923_out0 ? v_G1_2704_out0 : v_FF1_4721_out0;
always @(posedge clk) v_FF1_4722_out0 <= v_EN_2924_out0 ? v_G1_2705_out0 : v_FF1_4722_out0;
always @(posedge clk) v_FF1_4723_out0 <= v_EN_2925_out0 ? v_G1_2706_out0 : v_FF1_4723_out0;
always @(posedge clk) v_FF1_4724_out0 <= v_EN_2926_out0 ? v_G1_2707_out0 : v_FF1_4724_out0;
always @(posedge clk) v_FF1_4725_out0 <= v_EN_2927_out0 ? v_G1_2708_out0 : v_FF1_4725_out0;
always @(posedge clk) v_FF1_4726_out0 <= v_EN_2928_out0 ? v_G1_2709_out0 : v_FF1_4726_out0;
always @(posedge clk) v_FF1_4727_out0 <= v_EN_2929_out0 ? v_G1_2710_out0 : v_FF1_4727_out0;
always @(posedge clk) v_FF1_4728_out0 <= v_EN_2930_out0 ? v_G1_2711_out0 : v_FF1_4728_out0;
always @(posedge clk) v_FF1_4729_out0 <= v_EN_2931_out0 ? v_G1_2712_out0 : v_FF1_4729_out0;
always @(posedge clk) v_FF1_4730_out0 <= v_EN_2932_out0 ? v_G1_2713_out0 : v_FF1_4730_out0;
always @(posedge clk) v_FF1_4731_out0 <= v_EN_2933_out0 ? v_G1_2714_out0 : v_FF1_4731_out0;
always @(posedge clk) v_FF1_4732_out0 <= v_EN_2934_out0 ? v_G1_2715_out0 : v_FF1_4732_out0;
always @(posedge clk) v_REG3_4747_out0 <= v_D1_8842_out3 ? v_DIN3_10310_out0 : v_REG3_4747_out0;
always @(posedge clk) v_REG3_4748_out0 <= v_D1_8843_out3 ? v_DIN3_10311_out0 : v_REG3_4748_out0;
always @(posedge clk) v_FF7_4781_out0 <= v_ENABLE_2651_out0 ? v_MUX6_10976_out0 : v_FF7_4781_out0;
always @(posedge clk) v_FF1_4841_out0 <= v_G20_11040_out0;
always @(posedge clk) v_REG1_7031_out0 <= v_G8_7103_out0 ? v_MUX1_11061_out0 : v_REG1_7031_out0;
always @(posedge clk) v_FF5_7100_out0 <= v_ENABLE_2651_out0 ? v_MUX4_3219_out0 : v_FF5_7100_out0;
always @(posedge clk) v_REG1_7134_out0 <= v_EQ3_5861_out0 ? v_A1_11043_out0 : v_REG1_7134_out0;
always @(posedge clk) v_FF9_8805_out0 <= v_ENABLE_2651_out0 ? v_MUX8_2697_out0 : v_FF9_8805_out0;
always @(posedge clk) v_FF1_10325_out0 <= v_G3_2941_out0 ? v_G2_10799_out0 : v_FF1_10325_out0;
always @(posedge clk) v_FF1_10326_out0 <= v_G3_2942_out0 ? v_G2_10800_out0 : v_FF1_10326_out0;
always @(posedge clk) v_REG1_10368_out0 <= v__533_out0;
always @(posedge clk) v_REG1_10546_out0 <= v_G8_16_out0 ? v_OUT_3037_out0 : v_REG1_10546_out0;
always @(posedge clk) v_FF8_10849_out0 <= v_G21_3808_out0;
always @(posedge clk) v_FF8_10850_out0 <= v_G21_3809_out0;
always @(posedge clk) v_FF8_10851_out0 <= v_G21_3810_out0;
always @(posedge clk) v_FF8_10852_out0 <= v_G21_3811_out0;
always @(posedge clk) v_REG0_10912_out0 <= v_D1_8842_out0 ? v_DIN3_10310_out0 : v_REG0_10912_out0;
always @(posedge clk) v_REG0_10913_out0 <= v_D1_8843_out0 ? v_DIN3_10311_out0 : v_REG0_10913_out0;
always @(posedge clk) v_FF3_11046_out0 <= v_ENABLE_2651_out0 ? v_MUX2_4448_out0 : v_FF3_11046_out0;
always @(posedge clk) v_FF2_11062_out0 <= v_FF1_13511_out0;
always @(posedge clk) v_REG1_11130_out0 <= v_G2_6884_out0 ? v_COUT_3895_out0 : v_REG1_11130_out0;
always @(posedge clk) v_REG1_11131_out0 <= v_G2_6885_out0 ? v_COUT_3896_out0 : v_REG1_11131_out0;
always @(posedge clk) v_FF8_11222_out0 <= v_ENABLE_2651_out0 ? v_MUX7_10448_out0 : v_FF8_11222_out0;
always @(posedge clk) v_REG2_12251_out0 <= v_D1_8842_out2 ? v_DIN3_10310_out0 : v_REG2_12251_out0;
always @(posedge clk) v_REG2_12252_out0 <= v_D1_8843_out2 ? v_DIN3_10311_out0 : v_REG2_12252_out0;
always @(posedge clk) v_REG1_13338_out0 <= v_COUT_10922_out0;
always @(posedge clk) v_REG1_13339_out0 <= v_COUT_10937_out0;
v_RAM1_13398 I1 (v_RAM1_13398_out0, v_ADRESS_ins1_10617_out0, v_DATA_RAM_IN1_4779_out0, v_C3_2764_out0, clk);
always @(posedge clk) v_FF1_13511_out0 <= v_ROM1_462_out0;
assign v_C11_13766_out0 = 6'h0;
assign v_C11_13765_out0 = 6'h0;
assign v_C1_13447_out0 = 8'h0;
assign v_C1_13446_out0 = 8'h0;
assign v_C1_13278_out0 = 8'h0;
assign v_C1_13277_out0 = 8'h0;
assign v_C5_13267_out0 = 1'h1;
assign v_C1_11293_out0 = 2'h0;
assign v_C1_11292_out0 = 2'h0;
assign v_C10_11249_out0 = 5'h1f;
assign v_C10_11248_out0 = 5'h1f;
assign v_C2_11233_out0 = 3'h0;
assign v_C9_11160_out0 = 6'h3f;
assign v_C9_11159_out0 = 6'h3f;
assign v_C5_11031_out0 = 1'h0;
assign v_C3_10853_out0 = 3'h0;
assign v_C14_10796_out0 = 5'h1;
assign v_C14_10795_out0 = 5'h1;
assign v_C1_10790_out0 = 1'h0;
assign v_C1_10789_out0 = 1'h0;
assign v_C2_10762_out0 = 12'h7ff;
assign v_C2_10761_out0 = 12'h7ff;
assign v_C4_10619_out0 = 1'h1;
assign v_C5_10356_out0 = 2'h0;
assign v_C6_10318_out0 = 1'h1;
assign v_C6_10317_out0 = 1'h1;
assign v_C1_10316_out0 = 5'h0;
assign v_C1_10315_out0 = 5'h0;
assign v_C1_10314_out0 = 5'h0;
assign v_C1_10313_out0 = 5'h0;
assign v_C1_10306_out0 = 4'h0;
assign v_C1_10305_out0 = 4'h0;
assign v_C1_10267_out0 = 8'h0;
assign v_C1_10266_out0 = 8'h0;
assign v_C1_10259_out0 = 1'h0;
assign v_C1_8816_out0 = 1'h0;
assign v_C1_8815_out0 = 1'h0;
assign v_2_7072_out0 = 1'h1;
assign v_C1_6920_out0 = 4'h0;
assign v_C1_6919_out0 = 4'h0;
assign v_C1_6794_out0 = 2'h0;
assign v_C1_6793_out0 = 2'h0;
assign v_C3_4742_out0 = 1'h0;
assign v_C3_4741_out0 = 1'h0;
assign v_C11_4540_out0 = 16'hffff;
assign v_C11_4539_out0 = 16'hffff;
assign v_C7_3222_out0 = 1'h1;
assign v_C1_3211_out0 = 12'h0;
assign v_C1_3210_out0 = 12'h0;
assign v_C1_3206_out0 = 2'h0;
assign v_C1_3205_out0 = 2'h0;
assign v_C9_3030_out0 = 1'h0;
assign v_C9_3029_out0 = 1'h0;
assign v_C3_2764_out0 = 1'h0;
assign v_C8_2759_out0 = 5'h0;
assign v_C8_2758_out0 = 5'h0;
assign v_C1_2716_out0 = 3'h0;
assign v_C5_2689_out0 = 16'hffff;
assign v_C5_2688_out0 = 16'hffff;
assign v_C4_2594_out0 = 5'h0;
assign v_C4_2593_out0 = 5'h0;
assign v_C1_2427_out0 = 12'h7f4;
assign v_C1_2426_out0 = 12'h7f4;
assign v_C2_2413_out0 = 12'h0;
assign v_C7_2272_out0 = 1'h0;
assign v_C7_2271_out0 = 1'h0;
assign v_C13_2186_out0 = 16'h0;
assign v_C13_2185_out0 = 16'h0;
assign v_C12_2114_out0 = 6'hf;
assign v_C12_2113_out0 = 6'hf;
assign v_C1_2006_out0 = 4'h4;
assign v_C1_2005_out0 = 4'h4;
assign v_C7_1866_out0 = 16'h0;
assign v_C7_1865_out0 = 16'h0;
assign v_C10_1820_out0 = 1'h1;
assign v_C10_1819_out0 = 1'h1;
assign v_C_1808_out0 = 11'h0;
assign v_C_1807_out0 = 11'h0;
assign v_C6_1732_out0 = 1'h1;
assign v_C15_1731_out0 = 16'hffff;
assign v_C15_1730_out0 = 16'hffff;
assign v_C14_1675_out0 = 1'h1;
assign v_C14_1674_out0 = 1'h1;
assign v_C4_1201_out0 = 3'h0;
assign v_C12_1152_out0 = 1'h1;
assign v_C12_1151_out0 = 1'h1;
assign v_C1_607_out0 = 11'h0;
assign v_C1_606_out0 = 11'h0;
assign v_C1_605_out0 = 1'h0;
assign v_C1_604_out0 = 1'h0;
assign v_C1_436_out0 = 1'h1;
assign v_C13_406_out0 = 6'h31;
assign v_C13_405_out0 = 6'h31;
assign v_C4_90_out0 = 1'h0;
assign v_ROR_67_out0 = 2'h3;
assign v_ROR_66_out0 = 2'h3;
assign v_Q_291_out0 = v_FF1_4717_out0;
assign v_Q_292_out0 = v_FF1_4718_out0;
assign v_Q_293_out0 = v_FF1_4719_out0;
assign v_Q_294_out0 = v_FF1_4720_out0;
assign v_Q_295_out0 = v_FF1_4721_out0;
assign v_Q_296_out0 = v_FF1_4722_out0;
assign v_Q_297_out0 = v_FF1_4723_out0;
assign v_Q_298_out0 = v_FF1_4724_out0;
assign v_Q_299_out0 = v_FF1_4725_out0;
assign v_Q_300_out0 = v_FF1_4726_out0;
assign v_Q_301_out0 = v_FF1_4727_out0;
assign v_Q_302_out0 = v_FF1_4728_out0;
assign v_Q_303_out0 = v_FF1_4729_out0;
assign v_Q_304_out0 = v_FF1_4730_out0;
assign v_Q_305_out0 = v_FF1_4731_out0;
assign v_Q_306_out0 = v_FF1_4732_out0;
assign v_DATA_OUT_1135_out0 = v_data_ram_1818_out0;
assign v_EQ4_1142_out0 = v_REG1_7134_out0 == 12'h0;
assign v__1673_out0 = { v_FF1_4841_out0,v_C2_11233_out0 };
assign v_R0_1688_out0 = v_REG0_10912_out0;
assign v_R0_1689_out0 = v_REG0_10913_out0;
assign v_Q6_1889_out0 = v_FF7_2670_out0;
assign v_Q6_1890_out0 = v_FF7_2671_out0;
assign v_Q6_1891_out0 = v_FF7_2672_out0;
assign v_Q6_1892_out0 = v_FF7_2673_out0;
assign v_DIV_INST_2324_out0 = v_DIV_INST1_7011_out0;
assign v_DIV_INST_2325_out0 = v_DIV_INST0_6905_out0;
assign v_RAM_OUT1_2385_out0 = v_RAM1_13398_out0;
assign v_IR_2826_out0 = v_IHOLD_REGISTER_2013_out0;
assign v_IR_2827_out0 = v_IHOLD_REGISTER_2014_out0;
assign v__2887_out0 = { v_FF3_2016_out0,v_FF4_2106_out0 };
assign v__2888_out0 = { v_FF3_2017_out0,v_FF4_2107_out0 };
assign v__2959_out0 = v_REG1_2677_out0[0:0];
assign v__2959_out1 = v_REG1_2677_out0[7:7];
assign v_OUT_3037_out0 = v_REG1_2677_out0;
assign v_R2_3043_out0 = v_REG2_12251_out0;
assign v_R2_3044_out0 = v_REG2_12252_out0;
assign v_C_3197_out0 = v_REG1_11130_out0;
assign v_C_3198_out0 = v_REG1_11131_out0;
assign v_C_3207_out0 = v_REG1_11130_out0;
assign v_C_3208_out0 = v_REG1_11131_out0;
assign v_EQ1_3344_out0 = v_REG1_7031_out0 == 2'h2;
assign v_Q1_3993_out0 = v_FF1_4841_out0;
assign v_EN_4485_out0 = v_C5_13267_out0;
assign v_R3_4652_out0 = v_REG3_4747_out0;
assign v_R3_4653_out0 = v_REG3_4748_out0;
assign v_byte_ready_5842_out0 = v_C5_11031_out0;
assign v__5860_out0 = v_REG1_10368_out0[0:0];
assign v__5860_out1 = v_REG1_10368_out0[1:1];
assign v_Q7_6888_out0 = v_FF8_10849_out0;
assign v_Q7_6889_out0 = v_FF8_10850_out0;
assign v_Q7_6890_out0 = v_FF8_10851_out0;
assign v_Q7_6891_out0 = v_FF8_10852_out0;
assign v_NEG1_6921_out0 = v_C9_11159_out0;
assign v_NEG1_6922_out0 = v_C9_11160_out0;
assign v__7116_out0 = v_IHOLD_REGISTER_2013_out0[11:0];
assign v__7116_out1 = v_IHOLD_REGISTER_2013_out0[15:4];
assign v__7117_out0 = v_IHOLD_REGISTER_2014_out0[11:0];
assign v__7117_out1 = v_IHOLD_REGISTER_2014_out0[15:4];
assign v_RECEIVERSTREAM_7635_out0 = v_REG1_10546_out0;
assign v_RX_BYTEREADY_8756_out0 = v_FF1_4841_out0;
assign v_R1_8761_out0 = v_REG1_2314_out0;
assign v_R1_8762_out0 = v_REG1_2315_out0;
assign v_RAM_OUT0_8764_out0 = v_RAM0_1680_out0;
assign v_0B00001_10554_out0 = v_C14_10795_out0;
assign v_0B00001_10555_out0 = v_C14_10796_out0;
assign v_Q_10618_out0 = v_REG1_10368_out0;
assign v_0_10706_out0 = v_C7_2271_out0;
assign v_0_10707_out0 = v_C7_2272_out0;
assign v_G2_10799_out0 = ! v_FF1_10325_out0;
assign v_G2_10800_out0 = ! v_FF1_10326_out0;
assign {v_A1_11043_out1,v_A1_11043_out0 } = v_C2_2413_out0 + v_REG1_7134_out0 + v_C1_436_out0;
assign v_FLOAT_INST16_13443_out0 = v_FF1_10325_out0;
assign v_FLOAT_INST16_13444_out0 = v_FF1_10326_out0;
assign v_Q_13510_out0 = v_REG1_7031_out0;
assign v_STALL_DUAL_CORE_13618_out0 = v_C4_90_out0;
assign v_SEL2_280_out0 = v__7116_out0[9:9];
assign v_SEL2_281_out0 = v__7117_out0[9:9];
assign v_MEM_RAM_434_out0 = v_DATA_OUT_1135_out0;
assign v_MEM_RAM_435_out0 = v_DATA_OUT_1135_out0;
assign v_RECEIVER_STREAM_564_out0 = v_RECEIVERSTREAM_7635_out0;
assign v_Q_1153_out0 = v__2887_out0;
assign v_Q_1154_out0 = v__2888_out0;
assign v_G5_1198_out0 = ! v_EN_4485_out0;
assign v_Q2_1676_out0 = v_Q_291_out0;
assign v_Q2_1677_out0 = v_Q_295_out0;
assign v_Q2_1678_out0 = v_Q_299_out0;
assign v_Q2_1679_out0 = v_Q_303_out0;
assign v_G10_1943_out0 = !(v_Q_292_out0 || v_Q_291_out0);
assign v_G10_1944_out0 = !(v_Q_296_out0 || v_Q_295_out0);
assign v_G10_1945_out0 = !(v_Q_300_out0 || v_Q_299_out0);
assign v_G10_1946_out0 = !(v_Q_304_out0 || v_Q_303_out0);
assign v_G4_1960_out0 = v_Q_294_out0 && v_Q_292_out0;
assign v_G4_1961_out0 = v_Q_298_out0 && v_Q_296_out0;
assign v_G4_1962_out0 = v_Q_302_out0 && v_Q_300_out0;
assign v_G4_1963_out0 = v_Q_306_out0 && v_Q_304_out0;
assign v_G28_2098_out0 = v_Q7_6888_out0 && v_Q6_1889_out0;
assign v_G28_2099_out0 = v_Q7_6889_out0 && v_Q6_1890_out0;
assign v_G28_2100_out0 = v_Q7_6890_out0 && v_Q6_1891_out0;
assign v_G28_2101_out0 = v_Q7_6891_out0 && v_Q6_1892_out0;
assign v_RAM_OUT_2104_out0 = v_RAM_OUT1_2385_out0;
assign v_RAM_OUT_2105_out0 = v_RAM_OUT0_8764_out0;
assign v_Q1_2112_out0 = v__5860_out1;
assign v_EQ10_2320_out0 = v__7116_out1 == 4'h3;
assign v_EQ10_2321_out0 = v__7117_out1 == 4'h3;
assign v_RX_BYTE_READY_2436_out0 = v_RX_BYTEREADY_8756_out0;
assign v__2536_out0 = { v_EQ1_3344_out0,v_C1_2716_out0 };
assign v_COUT_2725_out0 = v_A1_11043_out1;
assign v_R3TEST_2872_out0 = v_R3_4652_out0;
assign v_R3TEST_2873_out0 = v_R3_4653_out0;
assign v_FLOAT_INST_2955_out0 = v_FLOAT_INST16_13443_out0;
assign v_FLOAT_INST_2956_out0 = v_FLOAT_INST16_13444_out0;
assign v_G2_2975_out0 = ((v_Q_294_out0 && !v_Q_292_out0) || (!v_Q_294_out0) && v_Q_292_out0);
assign v_G2_2976_out0 = ((v_Q_298_out0 && !v_Q_296_out0) || (!v_Q_298_out0) && v_Q_296_out0);
assign v_G2_2977_out0 = ((v_Q_302_out0 && !v_Q_300_out0) || (!v_Q_302_out0) && v_Q_300_out0);
assign v_G2_2978_out0 = ((v_Q_306_out0 && !v_Q_304_out0) || (!v_Q_306_out0) && v_Q_304_out0);
assign v__2983_out0 = v_Q_13510_out0[0:0];
assign v__2983_out1 = v_Q_13510_out0[1:1];
assign v_R0TEST_3184_out0 = v_R0_1688_out0;
assign v_R0TEST_3185_out0 = v_R0_1689_out0;
assign v_G2_4468_out0 = ! v_STALL_DUAL_CORE_13618_out0;
assign v_NOTUSED_4609_out0 = v__2959_out0;
assign v_EQ_4835_out0 = v__7116_out1 == 4'h0;
assign v_EQ_4836_out0 = v__7117_out1 == 4'h0;
assign v_G23_4852_out0 = ! v_Q7_6888_out0;
assign v_G23_4853_out0 = ! v_Q7_6889_out0;
assign v_G23_4854_out0 = ! v_Q7_6890_out0;
assign v_G23_4855_out0 = ! v_Q7_6891_out0;
assign v_RX_OVERFLOW_5848_out0 = v_EQ1_3344_out0;
assign v_EQ3_5861_out0 = v_Q_10618_out0 == 2'h3;
assign v_IR_7112_out0 = v_IR_2826_out0;
assign v_IR_7113_out0 = v_IR_2827_out0;
assign v__7183_out0 = { v_Q7_6888_out0,v_Q6_1889_out0 };
assign v__7184_out0 = { v_Q7_6889_out0,v_Q6_1890_out0 };
assign v__7185_out0 = { v_Q7_6890_out0,v_Q6_1891_out0 };
assign v__7186_out0 = { v_Q7_6891_out0,v_Q6_1892_out0 };
assign v_C_8648_out0 = v_C_3207_out0;
assign v_C_8649_out0 = v_C_3208_out0;
assign v_G1_8693_out0 = ! v_Q_294_out0;
assign v_G1_8694_out0 = ! v_Q_298_out0;
assign v_G1_8695_out0 = ! v_Q_302_out0;
assign v_G1_8696_out0 = ! v_Q_306_out0;
assign v_Q3_8737_out0 = v_Q_293_out0;
assign v_Q3_8738_out0 = v_Q_297_out0;
assign v_Q3_8739_out0 = v_Q_301_out0;
assign v_Q3_8740_out0 = v_Q_305_out0;
assign v_Q1_8859_out0 = v_Q_292_out0;
assign v_Q1_8860_out0 = v_Q_296_out0;
assign v_Q1_8861_out0 = v_Q_300_out0;
assign v_Q1_8862_out0 = v_Q_304_out0;
assign v_G9_10291_out0 = v_Q_294_out0 && v_Q_293_out0;
assign v_G9_10292_out0 = v_Q_298_out0 && v_Q_297_out0;
assign v_G9_10293_out0 = v_Q_302_out0 && v_Q_301_out0;
assign v_G9_10294_out0 = v_Q_306_out0 && v_Q_305_out0;
assign v_R1TEST_10485_out0 = v_R1_8761_out0;
assign v_R1TEST_10486_out0 = v_R1_8762_out0;
assign v_G24_10560_out0 = ((v_Q7_6888_out0 && !v_Q6_1889_out0) || (!v_Q7_6888_out0) && v_Q6_1889_out0);
assign v_G24_10561_out0 = ((v_Q7_6889_out0 && !v_Q6_1890_out0) || (!v_Q7_6889_out0) && v_Q6_1890_out0);
assign v_G24_10562_out0 = ((v_Q7_6890_out0 && !v_Q6_1891_out0) || (!v_Q7_6890_out0) && v_Q6_1891_out0);
assign v_G24_10563_out0 = ((v_Q7_6891_out0 && !v_Q6_1892_out0) || (!v_Q7_6891_out0) && v_Q6_1892_out0);
assign v_R2TEST_10708_out0 = v_R2_3043_out0;
assign v_R2TEST_10709_out0 = v_R2_3044_out0;
assign v_BYTE_READY_11172_out0 = v_byte_ready_5842_out0;
assign v_Q0_11198_out0 = v_Q_294_out0;
assign v_Q0_11199_out0 = v_Q_298_out0;
assign v_Q0_11200_out0 = v_Q_302_out0;
assign v_Q0_11201_out0 = v_Q_306_out0;
assign v_DIV_INSTRUCTION_11296_out0 = v_DIV_INST_2324_out0;
assign v_DIV_INSTRUCTION_11297_out0 = v_DIV_INST_2325_out0;
assign v_Q0_13351_out0 = v__5860_out0;
assign v_NOUSED_13492_out0 = v__7116_out0;
assign v_NOUSED_13493_out0 = v__7117_out0;
assign v_EQ2_8_out0 = v_Q_1153_out0 == 2'h2;
assign v_EQ2_9_out0 = v_Q_1154_out0 == 2'h2;
assign v_R3TEST_117_out0 = v_R3TEST_2872_out0;
assign v_R3TEST_118_out0 = v_R3TEST_2873_out0;
assign v_LS_204_out0 = v_EQ_4835_out0;
assign v_LS_205_out0 = v_EQ_4836_out0;
assign v_4BITCOUNTER_317_out0 = v__7183_out0;
assign v_4BITCOUNTER_318_out0 = v__7184_out0;
assign v_4BITCOUNTER_319_out0 = v__7185_out0;
assign v_4BITCOUNTER_320_out0 = v__7186_out0;
assign v_EQ4_611_out0 = v_Q_1153_out0 == 2'h0;
assign v_EQ4_612_out0 = v_Q_1154_out0 == 2'h0;
assign v_G6_1159_out0 = v_G4_1960_out0 && v_Q_291_out0;
assign v_G6_1160_out0 = v_G4_1961_out0 && v_Q_295_out0;
assign v_G6_1161_out0 = v_G4_1962_out0 && v_Q_299_out0;
assign v_G6_1162_out0 = v_G4_1963_out0 && v_Q_303_out0;
assign v_IR_1871_out0 = v_IR_7112_out0;
assign v_IR_1872_out0 = v_IR_7113_out0;
assign v_G12_2270_out0 = ! v_Q1_2112_out0;
assign v_EQ1_2540_out0 = v_Q_1153_out0 == 2'h1;
assign v_EQ1_2541_out0 = v_Q_1154_out0 == 2'h1;
assign v_STALL_DUAL_CORE_3128_out0 = v_G2_4468_out0;
assign v_G3_3343_out0 = v_G5_1198_out0 && v_Q1_2112_out0;
assign v_G38_3903_out0 = v_Q2_1676_out0 || v_Q3_8737_out0;
assign v_G38_3904_out0 = v_Q2_1677_out0 || v_Q3_8738_out0;
assign v_G38_3905_out0 = v_Q2_1678_out0 || v_Q3_8739_out0;
assign v_G38_3906_out0 = v_Q2_1679_out0 || v_Q3_8740_out0;
assign v_RX_OVERFLOW_4469_out0 = v_RX_OVERFLOW_5848_out0;
assign v_Q0_4470_out0 = v_Q0_11198_out0;
assign v_Q0_4471_out0 = v_Q0_11199_out0;
assign v_Q0_4472_out0 = v_Q0_11200_out0;
assign v_Q0_4473_out0 = v_Q0_11201_out0;
assign v_G6_4818_out0 = ! v__2983_out0;
assign v_C_4848_out0 = v_C_8648_out0;
assign v_C_4849_out0 = v_C_8649_out0;
assign v__5832_out0 = v_Q_1153_out0[0:0];
assign v__5832_out1 = v_Q_1153_out0[1:1];
assign v__5833_out0 = v_Q_1154_out0[0:0];
assign v__5833_out1 = v_Q_1154_out0[1:1];
assign v_Q2_6880_out0 = v_Q2_1676_out0;
assign v_Q2_6881_out0 = v_Q2_1677_out0;
assign v_Q2_6882_out0 = v_Q2_1678_out0;
assign v_Q2_6883_out0 = v_Q2_1679_out0;
assign v_G3_6894_out0 = ((v_G4_1960_out0 && !v_Q_291_out0) || (!v_G4_1960_out0) && v_Q_291_out0);
assign v_G3_6895_out0 = ((v_G4_1961_out0 && !v_Q_295_out0) || (!v_G4_1961_out0) && v_Q_295_out0);
assign v_G3_6896_out0 = ((v_G4_1962_out0 && !v_Q_299_out0) || (!v_G4_1962_out0) && v_Q_299_out0);
assign v_G3_6897_out0 = ((v_G4_1963_out0 && !v_Q_303_out0) || (!v_G4_1963_out0) && v_Q_303_out0);
assign v_G37_6900_out0 = v_Q1_8859_out0 || v_Q0_11198_out0;
assign v_G37_6901_out0 = v_Q1_8860_out0 || v_Q0_11199_out0;
assign v_G37_6902_out0 = v_Q1_8861_out0 || v_Q0_11200_out0;
assign v_G37_6903_out0 = v_Q1_8862_out0 || v_Q0_11201_out0;
assign v_Q1_6906_out0 = v_Q1_8859_out0;
assign v_Q1_6907_out0 = v_Q1_8860_out0;
assign v_Q1_6908_out0 = v_Q1_8861_out0;
assign v_Q1_6909_out0 = v_Q1_8862_out0;
assign v_G4_6914_out0 = ! v_Q0_13351_out0;
assign v_R0TEST_7005_out0 = v_R0TEST_3184_out0;
assign v_R0TEST_7006_out0 = v_R0TEST_3185_out0;
assign v_BYTE_READY_7021_out0 = v_BYTE_READY_11172_out0;
assign v_D_7680_out0 = v_G2_2975_out0;
assign v_D_7682_out0 = v_G1_8693_out0;
assign v_D_7684_out0 = v_G2_2976_out0;
assign v_D_7686_out0 = v_G1_8694_out0;
assign v_D_7688_out0 = v_G2_2977_out0;
assign v_D_7690_out0 = v_G1_8695_out0;
assign v_D_7692_out0 = v_G2_2978_out0;
assign v_D_7694_out0 = v_G1_8696_out0;
assign v_G11_8652_out0 = v_EN_4485_out0 && v_Q0_13351_out0;
assign v_G2_10278_out0 = ! v_EQ3_5861_out0;
assign v_RAM_OUT_10335_out0 = v_RAM_OUT_2104_out0;
assign v_RAM_OUT_10336_out0 = v_RAM_OUT_2105_out0;
assign v__10376_out0 = { v__1673_out0,v__2536_out0 };
assign v_FLOATING_INSTRUCTION_10391_out0 = v_FLOAT_INST_2955_out0;
assign v_FLOATING_INSTRUCTION_10392_out0 = v_FLOAT_INST_2956_out0;
assign v_EN_10451_out0 = v_G28_2098_out0;
assign v_EN_10452_out0 = v_G28_2099_out0;
assign v_EN_10453_out0 = v_G28_2100_out0;
assign v_EN_10454_out0 = v_G28_2101_out0;
assign v_G1_10476_out0 = ! v__2983_out1;
assign v_R1TEST_10498_out0 = v_R1TEST_10485_out0;
assign v_R1TEST_10499_out0 = v_R1TEST_10486_out0;
assign v_Q3_10518_out0 = v_Q3_8737_out0;
assign v_Q3_10519_out0 = v_Q3_8738_out0;
assign v_Q3_10520_out0 = v_Q3_8739_out0;
assign v_Q3_10521_out0 = v_Q3_8740_out0;
assign v_G8_10609_out0 = !(v_G9_10291_out0 && v_G10_1943_out0);
assign v_G8_10610_out0 = !(v_G9_10292_out0 && v_G10_1944_out0);
assign v_G8_10611_out0 = !(v_G9_10293_out0 && v_G10_1945_out0);
assign v_G8_10612_out0 = !(v_G9_10294_out0 && v_G10_1946_out0);
assign v_G8_10769_out0 = ! v_SEL2_280_out0;
assign v_G8_10770_out0 = ! v_SEL2_281_out0;
assign v_G1_10810_out0 = ((v_EN_4485_out0 && !v_Q0_13351_out0) || (!v_EN_4485_out0) && v_Q0_13351_out0);
assign v_G22_10983_out0 = v_G23_4852_out0 && v_Q6_1889_out0;
assign v_G22_10984_out0 = v_G23_4853_out0 && v_Q6_1890_out0;
assign v_G22_10985_out0 = v_G23_4854_out0 && v_Q6_1891_out0;
assign v_G22_10986_out0 = v_G23_4855_out0 && v_Q6_1892_out0;
assign v_R2TEST_10987_out0 = v_R2TEST_10708_out0;
assign v_R2TEST_10988_out0 = v_R2TEST_10709_out0;
assign v_RAM_OUT_11214_out0 = v_MEM_RAM_434_out0;
assign v_RAM_OUT_11215_out0 = v_MEM_RAM_435_out0;
assign v_BYTE_READY_13255_out0 = v_RX_BYTE_READY_2436_out0;
assign v_BYTE_RECEIVED_13441_out0 = v_RECEIVER_STREAM_564_out0;
assign v_SHIFHT_ENABLE_13500_out0 = v_G28_2098_out0;
assign v_SHIFHT_ENABLE_13501_out0 = v_G28_2099_out0;
assign v_SHIFHT_ENABLE_13502_out0 = v_G28_2100_out0;
assign v_SHIFHT_ENABLE_13503_out0 = v_G28_2101_out0;
assign v_EQ3_13504_out0 = v_Q_1153_out0 == 2'h3;
assign v_EQ3_13505_out0 = v_Q_1154_out0 == 2'h3;
assign v_DIV_INSTRUCTION_13635_out0 = v_DIV_INSTRUCTION_11296_out0;
assign v_DIV_INSTRUCTION_13636_out0 = v_DIV_INSTRUCTION_11297_out0;
assign v_EQ6_19_out0 = v_4BITCOUNTER_317_out0 == 2'h2;
assign v_R3_74_out0 = v_R3TEST_117_out0;
assign v_R3_75_out0 = v_R3TEST_118_out0;
assign v_NORMAL_181_out0 = v_EQ1_2540_out0;
assign v_NORMAL_182_out0 = v_EQ1_2541_out0;
assign v_LS_202_out0 = v_LS_204_out0;
assign v_LS_203_out0 = v_LS_205_out0;
assign v_Q1_307_out0 = v__5832_out1;
assign v_Q1_308_out0 = v__5833_out1;
assign v_RX_OVERFLOW_426_out0 = v_RX_OVERFLOW_4469_out0;
assign v_EXEC1LS_430_out0 = v_EQ2_8_out0;
assign v_EXEC1LS_431_out0 = v_EQ2_9_out0;
assign v_Q0_625_out0 = v__5832_out0;
assign v_Q0_626_out0 = v__5833_out0;
assign v_IR_640_out0 = v_IR_1871_out0;
assign v_IR_641_out0 = v_IR_1872_out0;
assign v_G7_1197_out0 = v_G11_8652_out0 && v_G12_2270_out0;
assign v_UNUSED3_1681_out0 = v_SHIFHT_ENABLE_13503_out0;
assign v_9_1700_out0 = v_G8_10609_out0;
assign v_9_1701_out0 = v_G8_10610_out0;
assign v_9_1702_out0 = v_G8_10611_out0;
assign v_9_1703_out0 = v_G8_10612_out0;
assign v_STALL_DUAL_CORE_1739_out0 = v_STALL_DUAL_CORE_3128_out0;
assign v_EQ9_2007_out0 = v_4BITCOUNTER_320_out0 == 2'h0;
assign v_R1_2056_out0 = v_R1TEST_10498_out0;
assign v_R1_2057_out0 = v_R1TEST_10499_out0;
assign v_G5_2584_out0 = ((v_G6_1159_out0 && !v_Q_293_out0) || (!v_G6_1159_out0) && v_Q_293_out0);
assign v_G5_2585_out0 = ((v_G6_1160_out0 && !v_Q_297_out0) || (!v_G6_1160_out0) && v_Q_297_out0);
assign v_G5_2586_out0 = ((v_G6_1161_out0 && !v_Q_301_out0) || (!v_G6_1161_out0) && v_Q_301_out0);
assign v_G5_2587_out0 = ((v_G6_1162_out0 && !v_Q_305_out0) || (!v_G6_1162_out0) && v_Q_305_out0);
assign v_R0_2850_out0 = v_R0TEST_7005_out0;
assign v_R0_2851_out0 = v_R0TEST_7006_out0;
assign v_G1_2911_out0 = v_EQ4_1142_out0 && v_G2_10278_out0;
assign v_EN_2919_out0 = v_EN_10451_out0;
assign v_EN_2920_out0 = v_EN_10451_out0;
assign v_EN_2921_out0 = v_EN_10451_out0;
assign v_EN_2922_out0 = v_EN_10451_out0;
assign v_EN_2923_out0 = v_EN_10452_out0;
assign v_EN_2924_out0 = v_EN_10452_out0;
assign v_EN_2925_out0 = v_EN_10452_out0;
assign v_EN_2926_out0 = v_EN_10452_out0;
assign v_EN_2927_out0 = v_EN_10453_out0;
assign v_EN_2928_out0 = v_EN_10453_out0;
assign v_EN_2929_out0 = v_EN_10453_out0;
assign v_EN_2930_out0 = v_EN_10453_out0;
assign v_EN_2931_out0 = v_EN_10454_out0;
assign v_EN_2932_out0 = v_EN_10454_out0;
assign v_EN_2933_out0 = v_EN_10454_out0;
assign v_EN_2934_out0 = v_EN_10454_out0;
assign v_START_3027_out0 = v_EQ4_611_out0;
assign v_START_3028_out0 = v_EQ4_612_out0;
assign v_RAM_OUT_3033_out0 = v_RAM_OUT_10335_out0;
assign v_RAM_OUT_3034_out0 = v_RAM_OUT_10336_out0;
assign v_G36_3135_out0 = !(v_G38_3903_out0 || v_G37_6900_out0);
assign v_G36_3136_out0 = !(v_G38_3904_out0 || v_G37_6901_out0);
assign v_G36_3137_out0 = !(v_G38_3905_out0 || v_G37_6902_out0);
assign v_G36_3138_out0 = !(v_G38_3906_out0 || v_G37_6903_out0);
assign v_EXEC2LS_3188_out0 = v_EQ3_13504_out0;
assign v_EXEC2LS_3189_out0 = v_EQ3_13505_out0;
assign v_UNUSED1_3220_out0 = v_SHIFHT_ENABLE_13502_out0;
assign v_EQ6_3257_out0 = v_4BITCOUNTER_319_out0 == 2'h0;
assign v_STALL_DUAL_CORE_3265_out0 = v_STALL_DUAL_CORE_3128_out0;
assign v_DIV_INSTRUCTION_3296_out0 = v_DIV_INSTRUCTION_13635_out0;
assign v_DIV_INSTRUCTION_3297_out0 = v_DIV_INSTRUCTION_13636_out0;
assign v_G7_6862_out0 = v_EQ_4835_out0 && v_G8_10769_out0;
assign v_G7_6863_out0 = v_EQ_4836_out0 && v_G8_10770_out0;
assign v_D_7679_out0 = v_G3_6894_out0;
assign v_D_7683_out0 = v_G3_6895_out0;
assign v_D_7687_out0 = v_G3_6896_out0;
assign v_D_7691_out0 = v_G3_6897_out0;
assign v_SHIFT_ENABLE_8684_out0 = v_SHIFHT_ENABLE_13500_out0;
assign v_EQ2_9795_out0 = v_4BITCOUNTER_317_out0 == 2'h1;
assign v__10287_out0 = { v_Q0_4470_out0,v_Q1_6906_out0 };
assign v__10288_out0 = { v_Q0_4471_out0,v_Q1_6907_out0 };
assign v__10289_out0 = { v_Q0_4472_out0,v_Q1_6908_out0 };
assign v__10290_out0 = { v_Q0_4473_out0,v_Q1_6909_out0 };
assign v_BYTE_READY_10558_out0 = v_BYTE_READY_7021_out0;
assign v_G10_10711_out0 = v_G4_6914_out0 && v_Q1_2112_out0;
assign v_R2_10904_out0 = v_R2TEST_10987_out0;
assign v_R2_10905_out0 = v_R2TEST_10988_out0;
assign v_EQ2_10981_out0 = v_4BITCOUNTER_318_out0 == 2'h0;
assign v_RESET_11174_out0 = v_G8_10609_out0;
assign v_RESET_11175_out0 = v_G8_10609_out0;
assign v_RESET_11176_out0 = v_G8_10609_out0;
assign v_RESET_11177_out0 = v_G8_10609_out0;
assign v_RESET_11178_out0 = v_G8_10610_out0;
assign v_RESET_11179_out0 = v_G8_10610_out0;
assign v_RESET_11180_out0 = v_G8_10610_out0;
assign v_RESET_11181_out0 = v_G8_10610_out0;
assign v_RESET_11182_out0 = v_G8_10611_out0;
assign v_RESET_11183_out0 = v_G8_10611_out0;
assign v_RESET_11184_out0 = v_G8_10611_out0;
assign v_RESET_11185_out0 = v_G8_10611_out0;
assign v_RESET_11186_out0 = v_G8_10612_out0;
assign v_RESET_11187_out0 = v_G8_10612_out0;
assign v_RESET_11188_out0 = v_G8_10612_out0;
assign v_RESET_11189_out0 = v_G8_10612_out0;
assign v_G9_13655_out0 = v_G6_4818_out0 && v__2983_out1;
assign v_BYTE_RECEIVED_13796_out0 = v_BYTE_RECEIVED_13441_out0;
assign v_FLOATING_INS_13797_out0 = v_FLOATING_INSTRUCTION_10391_out0;
assign v_FLOATING_INS_13798_out0 = v_FLOATING_INSTRUCTION_10392_out0;
assign v_R3_33_out0 = v_R3_74_out0;
assign v_R3_34_out0 = v_R3_75_out0;
assign v_MUX1_650_out0 = v_G1_2911_out0 ? v_C4_10619_out0 : v_FF2_11062_out0;
assign v_G1_1167_out0 = ! v_Q0_625_out0;
assign v_G1_1168_out0 = ! v_Q0_626_out0;
assign v_FLAOTING_INSTRUCTION_1859_out0 = v_FLOATING_INS_13797_out0;
assign v_FLAOTING_INSTRUCTION_1860_out0 = v_FLOATING_INS_13798_out0;
assign v_STALL_DUAL_CORE_1959_out0 = v_STALL_DUAL_CORE_1739_out0;
assign v_BYTE_RECEIVED_2231_out0 = v_BYTE_RECEIVED_13796_out0;
assign v_R0_2537_out0 = v_R0_2850_out0;
assign v_R0_2538_out0 = v_R0_2851_out0;
assign v_RAM_OUT_2628_out0 = v_RAM_OUT_3033_out0;
assign v_RAM_OUT_2629_out0 = v_RAM_OUT_3034_out0;
assign v_R1_2630_out0 = v_R1_2056_out0;
assign v_R1_2631_out0 = v_R1_2057_out0;
assign v_G1_2700_out0 = v_RESET_11174_out0 && v_D_7679_out0;
assign v_G1_2701_out0 = v_RESET_11175_out0 && v_D_7680_out0;
assign v_G1_2703_out0 = v_RESET_11177_out0 && v_D_7682_out0;
assign v_G1_2704_out0 = v_RESET_11178_out0 && v_D_7683_out0;
assign v_G1_2705_out0 = v_RESET_11179_out0 && v_D_7684_out0;
assign v_G1_2707_out0 = v_RESET_11181_out0 && v_D_7686_out0;
assign v_G1_2708_out0 = v_RESET_11182_out0 && v_D_7687_out0;
assign v_G1_2709_out0 = v_RESET_11183_out0 && v_D_7688_out0;
assign v_G1_2711_out0 = v_RESET_11185_out0 && v_D_7690_out0;
assign v_G1_2712_out0 = v_RESET_11186_out0 && v_D_7691_out0;
assign v_G1_2713_out0 = v_RESET_11187_out0 && v_D_7692_out0;
assign v_G1_2715_out0 = v_RESET_11189_out0 && v_D_7694_out0;
assign v_BYTE_READY_2852_out0 = v_BYTE_READY_10558_out0;
assign v_LS_2864_out0 = v_LS_202_out0;
assign v_LS_2865_out0 = v_LS_203_out0;
assign v_IR_2901_out0 = v_IR_640_out0;
assign v_IR_2902_out0 = v_IR_641_out0;
assign v__2960_out0 = { v__10287_out0,v_Q2_6880_out0 };
assign v__2961_out0 = { v__10288_out0,v_Q2_6881_out0 };
assign v__2962_out0 = { v__10289_out0,v_Q2_6882_out0 };
assign v__2963_out0 = { v__10290_out0,v_Q2_6883_out0 };
assign v_G6_4531_out0 = v_G10_10711_out0 || v_G3_3343_out0;
assign v_DIV_INSTRUCTION_4614_out0 = v_DIV_INSTRUCTION_3296_out0;
assign v_DIV_INSTRUCTION_4615_out0 = v_DIV_INSTRUCTION_3297_out0;
assign v_STALL_DUAL_CORE_4696_out0 = v_STALL_DUAL_CORE_1739_out0;
assign v_G2_6791_out0 = ! v_Q1_307_out0;
assign v_G2_6792_out0 = ! v_Q1_308_out0;
assign v_EXEC1LS_6795_out0 = v_EXEC1LS_430_out0;
assign v_EXEC1LS_6796_out0 = v_EXEC1LS_431_out0;
assign v_G13_7083_out0 = v_Q0_625_out0 && v_Q1_307_out0;
assign v_G13_7084_out0 = v_Q0_626_out0 && v_Q1_308_out0;
assign v_D_7681_out0 = v_G5_2584_out0;
assign v_D_7685_out0 = v_G5_2585_out0;
assign v_D_7689_out0 = v_G5_2586_out0;
assign v_D_7693_out0 = v_G5_2587_out0;
assign v_IR_7706_out0 = v_IR_640_out0;
assign v_IR_7707_out0 = v_IR_641_out0;
assign v_R2_10556_out0 = v_R2_10904_out0;
assign v_R2_10557_out0 = v_R2_10905_out0;
assign v_EXEC2LS_10979_out0 = v_EXEC2LS_3188_out0;
assign v_EXEC2LS_10980_out0 = v_EXEC2LS_3189_out0;
assign v_STALL_DUAL_CORE_12235_out0 = v_STALL_DUAL_CORE_3265_out0;
assign v_G9_13340_out0 = v_G7_6862_out0 && v_EXEC1LS_430_out0;
assign v_G9_13341_out0 = v_G7_6863_out0 && v_EXEC1LS_431_out0;
assign v_START_13394_out0 = v_START_3027_out0;
assign v_START_13395_out0 = v_START_3028_out0;
assign v_NORMAL_13429_out0 = v_NORMAL_181_out0;
assign v_NORMAL_13430_out0 = v_NORMAL_182_out0;
assign v_9_13623_out0 = v_9_1700_out0;
assign v_9_13624_out0 = v_9_1701_out0;
assign v_9_13625_out0 = v_9_1702_out0;
assign v_9_13626_out0 = v_9_1703_out0;
assign v__4_out0 = v_IR_2901_out0[14:12];
assign v__5_out0 = v_IR_2902_out0[14:12];
assign v_R3_27_out0 = v_R3_33_out0;
assign v_R3_28_out0 = v_R3_34_out0;
assign v_UNUSED_123_out0 = v_9_13625_out0;
assign v_G9_223_out0 = v_G6_4531_out0 || v_G7_1197_out0;
assign v_START_392_out0 = v_START_13394_out0;
assign v_START_393_out0 = v_START_13395_out0;
assign v_9_417_out0 = v_9_13624_out0;
assign v_LS_1202_out0 = v_LS_2864_out0;
assign v_LS_1203_out0 = v_LS_2865_out0;
assign v_G7_1684_out0 = v_G1_1167_out0 && v_Q1_307_out0;
assign v_G7_1685_out0 = v_G1_1168_out0 && v_Q1_308_out0;
assign v_G3_1720_out0 = ! v_FLAOTING_INSTRUCTION_1859_out0;
assign v_G3_1721_out0 = ! v_FLAOTING_INSTRUCTION_1860_out0;
assign v_R2_1726_out0 = v_R2_10556_out0;
assign v_R2_1727_out0 = v_R2_10557_out0;
assign v_RAM_OUT_1751_out0 = v_RAM_OUT_2628_out0;
assign v_RAM_OUT_1752_out0 = v_RAM_OUT_2629_out0;
assign v_UNUSED2_2424_out0 = v_9_13626_out0;
assign v__2599_out0 = v_IR_2901_out0[1:0];
assign v__2600_out0 = v_IR_2902_out0[1:0];
assign v_G1_2702_out0 = v_RESET_11176_out0 && v_D_7681_out0;
assign v_G1_2706_out0 = v_RESET_11180_out0 && v_D_7685_out0;
assign v_G1_2710_out0 = v_RESET_11184_out0 && v_D_7689_out0;
assign v_G1_2714_out0 = v_RESET_11188_out0 && v_D_7693_out0;
assign v_R1_2723_out0 = v_R1_2630_out0;
assign v_R1_2724_out0 = v_R1_2631_out0;
assign v__2773_out0 = { v__2960_out0,v_Q3_10518_out0 };
assign v__2774_out0 = { v__2961_out0,v_Q3_10519_out0 };
assign v__2775_out0 = { v__2962_out0,v_Q3_10520_out0 };
assign v__2776_out0 = { v__2963_out0,v_Q3_10521_out0 };
assign v_G2_3221_out0 = ! v_9_13623_out0;
assign v_EXEC2LS_3231_out0 = v_EXEC2LS_10979_out0;
assign v_EXEC2LS_3232_out0 = v_EXEC2LS_10980_out0;
assign v_wen_ram_4595_out0 = v_G9_13340_out0;
assign v_wen_ram_4596_out0 = v_G9_13341_out0;
assign v_IR1_6873_out0 = v_IR_7706_out0;
assign v_BIT_6918_out0 = v_MUX1_650_out0;
assign v_EXEC1_7029_out0 = v_EXEC1LS_6795_out0;
assign v_EXEC1_7030_out0 = v_EXEC1LS_6796_out0;
assign v__7095_out0 = v_IR_2901_out0[15:15];
assign v__7096_out0 = v_IR_2902_out0[15:15];
assign v_STALL_dual_core_8742_out0 = v_STALL_DUAL_CORE_1959_out0;
assign v_BYTE_RECEIVED_8819_out0 = v_BYTE_RECEIVED_2231_out0;
assign v_BYTE_RECEIVED_8820_out0 = v_BYTE_RECEIVED_2231_out0;
assign v_NORMAL_10256_out0 = v_NORMAL_13429_out0;
assign v_NORMAL_10257_out0 = v_NORMAL_13430_out0;
assign v__10371_out0 = { v_STALL_DUAL_CORE_4696_out0,v_C_1808_out0 };
assign v_EXEC1LS_10506_out0 = v_EXEC1LS_6795_out0;
assign v_EXEC1LS_10507_out0 = v_EXEC1LS_6796_out0;
assign v__10791_out0 = v_IR_2901_out0[11:10];
assign v__10792_out0 = v_IR_2902_out0[11:10];
assign v_G5_10914_out0 = v_Q0_625_out0 && v_G2_6791_out0;
assign v_G5_10915_out0 = v_Q0_626_out0 && v_G2_6792_out0;
assign v_BYTE_RECEIVED_11192_out0 = v_BYTE_RECEIVED_2231_out0;
assign v_STORE_12245_out0 = v_G9_13340_out0;
assign v_STORE_12246_out0 = v_G9_13341_out0;
assign v_R0_13295_out0 = v_R0_2537_out0;
assign v_R0_13296_out0 = v_R0_2538_out0;
assign v_IR0_13305_out0 = v_IR_7707_out0;
assign v_IR_13480_out0 = v_IR_2901_out0;
assign v_IR_13481_out0 = v_IR_2902_out0;
assign v_G3_13641_out0 = v_G1_1167_out0 && v_G2_6791_out0;
assign v_G3_13642_out0 = v_G1_1168_out0 && v_G2_6792_out0;
assign v_IR_105_out0 = v_IR_13480_out0;
assign v_IR_106_out0 = v_IR_13481_out0;
assign v__224_out0 = v_RAM_OUT_1751_out0[11:0];
assign v__224_out1 = v_RAM_OUT_1751_out0[15:4];
assign v__225_out0 = v_RAM_OUT_1752_out0[11:0];
assign v__225_out1 = v_RAM_OUT_1752_out0[15:4];
assign v_G1_277_out0 = v_EQ2_9795_out0 && v_G2_3221_out0;
assign v_R13_375_out0 = v_R3_27_out0;
assign v_R11_398_out0 = v_R1_2723_out0;
assign v__533_out0 = { v_G1_10810_out0,v_G9_223_out0 };
assign v_OP_621_out0 = v__4_out0;
assign v_OP_622_out0 = v__5_out0;
assign v_D_2108_out0 = v__10791_out0;
assign v_D_2109_out0 = v__10792_out0;
assign v_G16_2310_out0 = ! v_STORE_12245_out0;
assign v_G16_2311_out0 = ! v_STORE_12246_out0;
assign v__2422_out0 = v_IR_13480_out0[8:8];
assign v__2423_out0 = v_IR_13481_out0[8:8];
assign v_IR15_2464_out0 = v__7095_out0;
assign v_IR15_2465_out0 = v__7096_out0;
assign v_G8_2644_out0 = ! v_9_417_out0;
assign v__2846_out0 = v_IR_13480_out0[4:0];
assign v__2847_out0 = v_IR_13481_out0[4:0];
assign v_G6_2905_out0 = v_G3_13641_out0 || v_G7_1684_out0;
assign v_G6_2906_out0 = v_G3_13642_out0 || v_G7_1685_out0;
assign v_LS1_3169_out0 = v_LS_1202_out0;
assign v_BIT_IN1_3209_out0 = v_BIT_6918_out0;
assign v_NORMAL_3353_out0 = v_NORMAL_10256_out0;
assign v_NORMAL_3354_out0 = v_NORMAL_10257_out0;
assign v_R00_3807_out0 = v_R0_13296_out0;
assign v__3942_out0 = v_IR_13480_out0[7:4];
assign v__3943_out0 = v_IR_13481_out0[7:4];
assign v_LS0_4548_out0 = v_LS_1203_out0;
assign v__4837_out0 = v_IR_13480_out0[9:9];
assign v__4838_out0 = v_IR_13481_out0[9:9];
assign v_SEL1_5798_out0 = v_IR_13480_out0[15:12];
assign v_SEL1_5799_out0 = v_IR_13481_out0[15:12];
assign v_R02_6966_out0 = v_R2_1727_out0;
assign v_WEN_RAM_7079_out0 = v_wen_ram_4595_out0;
assign v_WEN_RAM_7080_out0 = v_wen_ram_4596_out0;
assign v_EN_7094_out0 = v_STALL_dual_core_8742_out0;
assign v_BYTE_RECEIVED_7101_out0 = v_BYTE_RECEIVED_8819_out0;
assign v_BYTE_RECEIVED_7102_out0 = v_BYTE_RECEIVED_8820_out0;
assign v_M_7177_out0 = v__2599_out0;
assign v_M_7178_out0 = v__2600_out0;
assign v_R12_10714_out0 = v_R2_1726_out0;
assign v_EXEC1_10763_out0 = v_EXEC1_7029_out0;
assign v_EXEC1_10764_out0 = v_EXEC1_7030_out0;
assign v_A_10822_out0 = v__10371_out0;
assign v_EXEC1LS_10843_out0 = v_EXEC1LS_10506_out0;
assign v_EXEC1LS_10844_out0 = v_EXEC1LS_10507_out0;
assign v__11163_out0 = v_IR_13480_out0[3:2];
assign v__11164_out0 = v_IR_13481_out0[3:2];
assign v_R10_11216_out0 = v_R0_13295_out0;
assign v_8BITCOUNTER_13281_out0 = v__2773_out0;
assign v_8BITCOUNTER_13282_out0 = v__2774_out0;
assign v_8BITCOUNTER_13283_out0 = v__2775_out0;
assign v_8BITCOUNTER_13284_out0 = v__2776_out0;
assign v_R03_13304_out0 = v_R3_28_out0;
assign v_EXEC2LS_13558_out0 = v_EXEC2LS_3231_out0;
assign v_EXEC2LS_13559_out0 = v_EXEC2LS_3232_out0;
assign v_WRITE_EN_13653_out0 = v_wen_ram_4595_out0;
assign v_WRITE_EN_13654_out0 = v_wen_ram_4596_out0;
assign v_R01_13752_out0 = v_R1_2724_out0;
assign v__61_out0 = v_A_10822_out0[10:10];
assign v__172_out0 = v_A_10822_out0[7:7];
assign v__180_out0 = v_A_10822_out0[3:3];
assign v_B_273_out0 = v__3942_out0;
assign v_B_274_out0 = v__3943_out0;
assign v__288_out0 = v_A_10822_out0[2:2];
assign v_EQ1_315_out0 = v__224_out1 == 4'h0;
assign v_EQ1_316_out0 = v__225_out1 == 4'h0;
assign v_G15_1855_out0 = !(v_EXEC1_10763_out0 || v_FF1_48_out0);
assign v_G15_1856_out0 = !(v_EXEC1_10764_out0 || v_FF1_49_out0);
assign v_EQ1_1857_out0 = v_SEL1_5798_out0 == 4'h1;
assign v_EQ1_1858_out0 = v_SEL1_5799_out0 == 4'h1;
assign v__1876_out0 = v_A_10822_out0[11:11];
assign v_EQ6_1966_out0 = v__224_out1 == 4'h5;
assign v_EQ6_1967_out0 = v__225_out1 == 4'h5;
assign v__2023_out0 = v_A_10822_out0[5:5];
assign v_EXEC2_2110_out0 = v_EXEC2LS_13558_out0;
assign v_EXEC2_2111_out0 = v_EXEC2LS_13559_out0;
assign v_EQ4_2149_out0 = v_8BITCOUNTER_13281_out0 == 4'h0;
assign v__2269_out0 = v_A_10822_out0[8:8];
assign v_EQ9_2390_out0 = v__224_out1 == 4'h3;
assign v_EQ9_2391_out0 = v__225_out1 == 4'h3;
assign v_EQ8_2453_out0 = v__224_out1 == 4'h7;
assign v_EQ8_2454_out0 = v__225_out1 == 4'h7;
assign v_EQ11_2456_out0 = v__224_out1 == 4'h1;
assign v_EQ11_2457_out0 = v__225_out1 == 4'h1;
assign v_IN_2466_out0 = v_BIT_IN1_3209_out0;
assign v_ADRESS_2542_out0 = v__224_out0;
assign v_ADRESS_2543_out0 = v__225_out0;
assign v_G21_2656_out0 = ! v_WEN_RAM_7079_out0;
assign v_G21_2657_out0 = ! v_WEN_RAM_7080_out0;
assign v_WEN_2765_out0 = v_WRITE_EN_13653_out0;
assign v_WEN_2766_out0 = v_WRITE_EN_13654_out0;
assign v_EXEC2LS_2844_out0 = v_EXEC2LS_13558_out0;
assign v_EXEC2LS_2845_out0 = v_EXEC2LS_13559_out0;
assign v_EQ8_2874_out0 = v_8BITCOUNTER_13284_out0 == 4'h0;
assign v_SEL1_2914_out0 = v__224_out0[9:9];
assign v_SEL1_2915_out0 = v__225_out0[9:9];
assign v_EQ3_2966_out0 = v_SEL1_5798_out0 == 4'h9;
assign v_EQ3_2967_out0 = v_SEL1_5799_out0 == 4'h9;
assign v__3124_out0 = v_A_10822_out0[1:1];
assign v_EXEC2_3170_out0 = v_NORMAL_3353_out0;
assign v_EXEC2_3171_out0 = v_NORMAL_3354_out0;
assign v_EQ4_3227_out0 = v_SEL1_5798_out0 == 4'h8;
assign v_EQ4_3228_out0 = v_SEL1_5799_out0 == 4'h8;
assign v__3271_out0 = v_A_10822_out0[4:4];
assign v_EQ7_3307_out0 = v__224_out1 == 4'h6;
assign v_EQ7_3308_out0 = v__225_out1 == 4'h6;
assign v_exec1ls_3341_out0 = v_EXEC1LS_10843_out0;
assign v_exec1ls_3342_out0 = v_EXEC1LS_10844_out0;
assign v_EXEC1LS_4697_out0 = v_EXEC1LS_10843_out0;
assign v_EXEC1LS_4698_out0 = v_EXEC1LS_10844_out0;
assign v_EQ5_4860_out0 = v__224_out1 == 4'h4;
assign v_EQ5_4861_out0 = v__225_out1 == 4'h4;
assign v_K_5792_out0 = v__2846_out0;
assign v_K_5793_out0 = v__2847_out0;
assign v__7081_out0 = { v_BYTE_RECEIVED_7101_out0,v_C1_13277_out0 };
assign v__7082_out0 = { v_BYTE_RECEIVED_7102_out0,v_C1_13278_out0 };
assign v_NORMAL_7114_out0 = v_NORMAL_3353_out0;
assign v_NORMAL_7115_out0 = v_NORMAL_3354_out0;
assign v_EXEC1_7128_out0 = v_EXEC1LS_10843_out0;
assign v_EXEC1_7129_out0 = v_EXEC1LS_10844_out0;
assign v_EQ3_7145_out0 = v__224_out1 == 4'h2;
assign v_EQ3_7146_out0 = v__225_out1 == 4'h2;
assign v_C_8653_out0 = v__4837_out0;
assign v_C_8654_out0 = v__4838_out0;
assign v_SHIFT_8661_out0 = v__11163_out0;
assign v_SHIFT_8662_out0 = v__11164_out0;
assign v_D_8752_out0 = v_D_2108_out0;
assign v_D_8753_out0 = v_D_2109_out0;
assign v__9791_out0 = { v_C1_13277_out0,v_BYTE_RECEIVED_7101_out0 };
assign v__9792_out0 = { v_C1_13278_out0,v_BYTE_RECEIVED_7102_out0 };
assign v_EQ1_10329_out0 = v_8BITCOUNTER_13282_out0 == 4'h0;
assign v_LDR_STR0_10349_out0 = v_LS0_4548_out0;
assign v_AD2_10699_out0 = v_M_7177_out0;
assign v_AD2_10700_out0 = v_M_7178_out0;
assign v_IR_10816_out0 = v_IR_105_out0;
assign v_IR_10817_out0 = v_IR_106_out0;
assign v_OP_11223_out0 = v_OP_621_out0;
assign v_OP_11224_out0 = v_OP_622_out0;
assign v__11243_out0 = v_A_10822_out0[9:9];
assign v_S_11300_out0 = v__2422_out0;
assign v_S_11301_out0 = v__2423_out0;
assign v__13397_out0 = v_A_10822_out0[6:6];
assign v__13563_out0 = v_A_10822_out0[0:0];
assign v_LDR_STR1_13616_out0 = v_LS1_3169_out0;
assign v_EQ7_13769_out0 = v_8BITCOUNTER_13283_out0 == 4'h0;
assign v_AD1_13774_out0 = v_D_2108_out0;
assign v_AD1_13775_out0 = v_D_2109_out0;
assign v_BIT_STREAM_IN_13_out0 = v_IN_2466_out0;
assign v_G4_381_out0 = v_EQ3_2966_out0 || v_EQ4_3227_out0;
assign v_G4_382_out0 = v_EQ3_2967_out0 || v_EQ4_3228_out0;
assign v_G20_598_out0 = v_EXEC1_10763_out0 && v_G21_2656_out0;
assign v_G20_599_out0 = v_EXEC1_10764_out0 && v_G21_2657_out0;
assign v_EXEC20_629_out0 = v_EXEC2_2111_out0;
assign v_B_1155_out0 = v_B_273_out0;
assign v_B_1156_out0 = v_B_274_out0;
assign v_EQ6_1686_out0 = v_OP_11223_out0 == 3'h5;
assign v_EQ6_1687_out0 = v_OP_11224_out0 == 3'h5;
assign v__1724_out0 = v_IR_10816_out0[14:14];
assign v__1725_out0 = v_IR_10817_out0[14:14];
assign v_JMI_1939_out0 = v_EQ6_1966_out0;
assign v_JMI_1940_out0 = v_EQ6_1967_out0;
assign v_EXEC2_2010_out0 = v_EXEC2_3170_out0;
assign v_EXEC2_2011_out0 = v_EXEC2_3171_out0;
assign v_NORMAL0_2307_out0 = v_NORMAL_7115_out0;
assign v_EXEC10_2329_out0 = v_exec1ls_3342_out0;
assign v_ADRESS_2339_out0 = v_ADRESS_2542_out0;
assign v_ADRESS_2340_out0 = v_ADRESS_2543_out0;
assign v__2430_out0 = v_IR_10816_out0[15:15];
assign v__2431_out0 = v_IR_10817_out0[15:15];
assign v__2470_out0 = v_IR_10816_out0[13:13];
assign v__2471_out0 = v_IR_10817_out0[13:13];
assign v_K_2636_out0 = v_K_5792_out0;
assign v_K_2637_out0 = v_K_5793_out0;
assign v_G2_2652_out0 = v_EQ9_2390_out0 || v_EQ10_2320_out0;
assign v_G2_2653_out0 = v_EQ9_2391_out0 || v_EQ10_2321_out0;
assign v_SUB_2695_out0 = v_EQ3_2966_out0;
assign v_SUB_2696_out0 = v_EQ3_2967_out0;
assign v_G5_2756_out0 = ! v_SEL1_2914_out0;
assign v_G5_2757_out0 = ! v_SEL1_2915_out0;
assign v__2831_out0 = v_AD2_10699_out0[0:0];
assign v__2831_out1 = v_AD2_10699_out0[1:1];
assign v__2832_out0 = v_AD2_10700_out0[0:0];
assign v__2832_out1 = v_AD2_10700_out0[1:1];
assign v__2860_out0 = v_IR_10816_out0[12:12];
assign v__2861_out0 = v_IR_10817_out0[12:12];
assign v_EQ8_2951_out0 = v_OP_11223_out0 == 3'h7;
assign v_EQ8_2952_out0 = v_OP_11224_out0 == 3'h7;
assign v_MULTI_OPCODE_3020_out0 = v_EQ1_1857_out0;
assign v_MULTI_OPCODE_3021_out0 = v_EQ1_1858_out0;
assign v_EXEC1_3038_out0 = v_EXEC1_7128_out0;
assign v_EXEC1_3039_out0 = v_EXEC1_7129_out0;
assign v_EXEC2LS_3081_out0 = v_EXEC2LS_2844_out0;
assign v_EXEC2LS_3082_out0 = v_EXEC2LS_2845_out0;
assign v__3897_out0 = v_IR_10816_out0[9:0];
assign v__3897_out1 = v_IR_10816_out0[15:6];
assign v__3898_out0 = v_IR_10817_out0[9:0];
assign v__3898_out1 = v_IR_10817_out0[15:6];
assign v_EXEC11_4528_out0 = v_exec1ls_3341_out0;
assign v_FLOAT_4603_out0 = v_EQ3_7145_out0;
assign v_FLOAT_4604_out0 = v_EQ3_7146_out0;
assign v_G25_4658_out0 = v_EQ8_2874_out0 && v_EQ9_2007_out0;
assign v_NORMAL1_6790_out0 = v_NORMAL_7114_out0;
assign v_REN1_6874_out0 = v_LDR_STR1_13616_out0;
assign v__6876_out0 = v_AD1_13774_out0[0:0];
assign v__6876_out1 = v_AD1_13774_out0[1:1];
assign v__6877_out0 = v_AD1_13775_out0[0:0];
assign v__6877_out1 = v_AD1_13775_out0[1:1];
assign v_EQ1_7098_out0 = v_OP_11223_out0 == 3'h0;
assign v_EQ1_7099_out0 = v_OP_11224_out0 == 3'h0;
assign v_EQ3_7126_out0 = v_OP_11223_out0 == 3'h2;
assign v_EQ3_7127_out0 = v_OP_11224_out0 == 3'h2;
assign v_JMP_8825_out0 = v_EQ5_4860_out0;
assign v_JMP_8826_out0 = v_EQ5_4861_out0;
assign v_EQ4_10345_out0 = v_OP_11223_out0 == 3'h3;
assign v_EQ4_10346_out0 = v_OP_11224_out0 == 3'h3;
assign v_STP_10352_out0 = v_EQ8_2453_out0;
assign v_STP_10353_out0 = v_EQ8_2454_out0;
assign v_EQ5_10364_out0 = v_OP_11223_out0 == 3'h4;
assign v_EQ5_10365_out0 = v_OP_11224_out0 == 3'h4;
assign v_EQ7_10399_out0 = v_OP_11223_out0 == 3'h6;
assign v_EQ7_10400_out0 = v_OP_11224_out0 == 3'h6;
assign v_JEQ_10496_out0 = v_EQ7_3307_out0;
assign v_JEQ_10497_out0 = v_EQ7_3308_out0;
assign v_RD_10522_out0 = v_D_8752_out0;
assign v_RD_10523_out0 = v_D_8753_out0;
assign v_EXEC2LS_10549_out0 = v_EXEC2_2110_out0;
assign v_SHIFT_10615_out0 = v_SHIFT_8661_out0;
assign v_SHIFT_10616_out0 = v_SHIFT_8662_out0;
assign v_G22_10620_out0 = v_EQ7_13769_out0 && v_EQ6_3257_out0;
assign v_EXEC1LS_10703_out0 = v_EXEC1LS_4697_out0;
assign v_EXEC1LS_10704_out0 = v_EXEC1LS_4698_out0;
assign v_EQ2_10771_out0 = v_OP_11223_out0 == 3'h1;
assign v_EQ2_10772_out0 = v_OP_11224_out0 == 3'h1;
assign v_G5_10989_out0 = ! v_EQ4_2149_out0;
assign v_WEN_11038_out0 = v_WEN_2765_out0;
assign v_WEN_11039_out0 = v_WEN_2766_out0;
assign v_REN0_11136_out0 = v_LDR_STR0_10349_out0;
assign v_G1_11157_out0 = v_EQ1_315_out0 || v_EQ9_2390_out0;
assign v_G1_11158_out0 = v_EQ1_316_out0 || v_EQ9_2391_out0;
assign v_G9_13564_out0 = v_EQ2_10981_out0 && v_EQ1_10329_out0;
assign v_C_13767_out0 = v_C_8653_out0;
assign v_C_13768_out0 = v_C_8654_out0;
assign v_G8_16_out0 = v_G1_277_out0 && v_BIT_STREAM_IN_13_out0;
assign v_STP_52_out0 = v_STP_10352_out0;
assign v_STP_53_out0 = v_STP_10353_out0;
assign v__124_out0 = { v_K_2636_out0,v_C1_606_out0 };
assign v__125_out0 = { v_K_2637_out0,v_C1_607_out0 };
assign v_C_238_out0 = v_C_13767_out0;
assign v_C_239_out0 = v_C_13768_out0;
assign v_MUX4_376_out0 = v__2831_out0 ? v_R1_8761_out0 : v_R0_1688_out0;
assign v_MUX4_377_out0 = v__2832_out0 ? v_R1_8762_out0 : v_R0_1689_out0;
assign v_EXEC2_441_out0 = v_EXEC2_2010_out0;
assign v_EXEC2_442_out0 = v_EXEC2_2011_out0;
assign v_G4_1667_out0 = v_EQ1_315_out0 && v_G5_2756_out0;
assign v_G4_1668_out0 = v_EQ1_316_out0 && v_G5_2757_out0;
assign v_UART_1823_out0 = v_G2_2652_out0;
assign v_UART_1824_out0 = v_G2_2653_out0;
assign v_EXEC1_1863_out0 = v_EXEC1LS_10703_out0;
assign v_EXEC1_1864_out0 = v_EXEC1LS_10704_out0;
assign v_G3_1949_out0 = v_EQ11_2456_out0 || v_G1_11157_out0;
assign v_G3_1950_out0 = v_EQ11_2457_out0 || v_G1_11158_out0;
assign v_JEQ_2234_out0 = v_JEQ_10496_out0;
assign v_JEQ_2235_out0 = v_JEQ_10497_out0;
assign v_BIT_2328_out0 = v_BIT_STREAM_IN_13_out0;
assign v_G7_2455_out0 = v_G9_13564_out0 || v_G8_2644_out0;
assign v_MUX1_2532_out0 = v__6876_out0 ? v_REG1_2314_out0 : v_REG0_10912_out0;
assign v_MUX1_2533_out0 = v__6877_out0 ? v_REG1_2315_out0 : v_REG0_10913_out0;
assign v_WEN0_2588_out0 = v_WEN_11039_out0;
assign v_EXEC1_2634_out0 = v_EXEC1LS_10703_out0;
assign v_EXEC1_2635_out0 = v_EXEC1LS_10704_out0;
assign v_EXEC2_2647_out0 = v_EXEC2LS_3081_out0;
assign v_EXEC2_2648_out0 = v_EXEC2LS_3082_out0;
assign v_NOTUSED_2698_out0 = v__3897_out1;
assign v_NOTUSED_2699_out0 = v__3898_out1;
assign v_SUB_INSTRUCTION_2789_out0 = v_SUB_2695_out0;
assign v_SUB_INSTRUCTION_2790_out0 = v_SUB_2696_out0;
assign v_EXEC11_2830_out0 = v_EXEC11_4528_out0;
assign v_JMP_3233_out0 = v_JMP_8825_out0;
assign v_JMP_3234_out0 = v_JMP_8826_out0;
assign v_EXEC2_3241_out0 = v_EXEC2LS_3081_out0;
assign v_EXEC2_3242_out0 = v_EXEC2LS_3082_out0;
assign v_TST_3819_out0 = v_EQ8_2951_out0;
assign v_TST_3820_out0 = v_EQ8_2952_out0;
assign v_AND_3858_out0 = v_EQ7_10399_out0;
assign v_AND_3859_out0 = v_EQ7_10400_out0;
assign v_MULTI_INSTRUCTION_3953_out0 = v_MULTI_OPCODE_3020_out0;
assign v_MULTI_INSTRUCTION_3954_out0 = v_MULTI_OPCODE_3021_out0;
assign v_G24_3955_out0 = ! v__2470_out0;
assign v_G24_3956_out0 = ! v__2471_out0;
assign v_G3_3959_out0 = v_G4_381_out0 && v_FLOATING_INS_13797_out0;
assign v_G3_3960_out0 = v_G4_382_out0 && v_FLOATING_INS_13798_out0;
assign v_ADD_4455_out0 = v_EQ1_7098_out0;
assign v_ADD_4456_out0 = v_EQ1_7099_out0;
assign v__4526_out0 = v__3897_out0[8:0];
assign v__4526_out1 = v__3897_out0[9:1];
assign v__4527_out0 = v__3898_out0[8:0];
assign v__4527_out1 = v__3898_out0[9:1];
assign v_MUX2_4612_out0 = v__6876_out0 ? v_REG3_4747_out0 : v_REG2_12251_out0;
assign v_MUX2_4613_out0 = v__6877_out0 ? v_REG3_4748_out0 : v_REG2_12252_out0;
assign v_BIN_5853_out0 = v_B_1155_out0;
assign v_BIN_5854_out0 = v_B_1156_out0;
assign v_G28_6868_out0 = ! v__1724_out0;
assign v_G28_6869_out0 = ! v__1725_out0;
assign v_G25_6962_out0 = v__2430_out0 && v__1724_out0;
assign v_G25_6963_out0 = v__2431_out0 && v__1725_out0;
assign v_JUMPADRESS_6964_out0 = v_ADRESS_2339_out0;
assign v_JUMPADRESS_6965_out0 = v_ADRESS_2340_out0;
assign v_STARTBIT_6967_out0 = v_BIT_STREAM_IN_13_out0;
assign v_FLOAT_7676_out0 = v_FLOAT_4603_out0;
assign v_FLOAT_7677_out0 = v_FLOAT_4604_out0;
assign v_SUB_8663_out0 = v_EQ2_10771_out0;
assign v_SUB_8664_out0 = v_EQ2_10772_out0;
assign v_WEN1_8763_out0 = v_WEN_11038_out0;
assign v_EXEC10_8812_out0 = v_EXEC10_2329_out0;
assign v_MUX5_8840_out0 = v__2831_out0 ? v_R3_4652_out0 : v_R2_3043_out0;
assign v_MUX5_8841_out0 = v__2832_out0 ? v_R3_4653_out0 : v_R2_3044_out0;
assign v_MOV_10389_out0 = v_EQ5_10364_out0;
assign v_MOV_10390_out0 = v_EQ5_10365_out0;
assign v_ADC_10393_out0 = v_EQ3_7126_out0;
assign v_ADC_10394_out0 = v_EQ3_7127_out0;
assign v_G3_10462_out0 = v_G5_10989_out0 && v_EQ6_19_out0;
assign v_G21_10681_out0 = ! v_G22_10620_out0;
assign v_MULTI_OPCODE_11096_out0 = v_MULTI_OPCODE_3020_out0;
assign v_MULTI_OPCODE_11097_out0 = v_MULTI_OPCODE_3021_out0;
assign v_G2_12230_out0 = v_EXEC2_2010_out0 || v_EXEC2LS_3081_out0;
assign v_G2_12231_out0 = v_EXEC2_2011_out0 || v_EXEC2LS_3082_out0;
assign v_JMI_13349_out0 = v_JMI_1939_out0;
assign v_JMI_13350_out0 = v_JMI_1940_out0;
assign v_SBC_13605_out0 = v_EQ4_10345_out0;
assign v_SBC_13606_out0 = v_EQ4_10346_out0;
assign v_CMP_13609_out0 = v_EQ6_1686_out0;
assign v_CMP_13610_out0 = v_EQ6_1687_out0;
assign v_EXEC1_20_out0 = v_EXEC1_1863_out0;
assign v_EXEC1_21_out0 = v_EXEC1_1864_out0;
assign v_JMI_88_out0 = v_JMI_13349_out0;
assign v_JMI_89_out0 = v_JMI_13350_out0;
assign v_MOV_196_out0 = v_MOV_10389_out0;
assign v_MOV_197_out0 = v_MOV_10390_out0;
assign v_MUX3_313_out0 = v__6876_out1 ? v_MUX2_4612_out0 : v_MUX1_2532_out0;
assign v_MUX3_314_out0 = v__6877_out1 ? v_MUX2_4613_out0 : v_MUX1_2533_out0;
assign v_C_379_out0 = v_C_238_out0;
assign v_C_380_out0 = v_C_239_out0;
assign v_STALL_427_out0 = v_G3_1949_out0;
assign v_STALL_428_out0 = v_G3_1950_out0;
assign v_MUX1_534_out0 = v_C_238_out0 ? v_ROR_66_out0 : v_SHIFT_10615_out0;
assign v_MUX1_535_out0 = v_C_239_out0 ? v_ROR_67_out0 : v_SHIFT_10616_out0;
assign v_JMP_546_out0 = v_JMP_3233_out0;
assign v_JMP_547_out0 = v_JMP_3234_out0;
assign v_G18_567_out0 = v_EXEC11_2830_out0 && v_REN1_6874_out0;
assign v_FLOATING_EN_ALU_634_out0 = v_G3_3959_out0;
assign v_FLOATING_EN_ALU_635_out0 = v_G3_3960_out0;
assign v_MUX2_1145_out0 = v_G2_12230_out0 ? v_D_2108_out0 : v_M_7177_out0;
assign v_MUX2_1146_out0 = v_G2_12231_out0 ? v_D_2109_out0 : v_M_7178_out0;
assign v_EQ1_1157_out0 = v__4526_out1 == 1'h0;
assign v_EQ1_1158_out0 = v__4527_out1 == 1'h0;
assign v_G1_2225_out0 = ! v_TST_3819_out0;
assign v_G1_2226_out0 = ! v_TST_3820_out0;
assign v_MUX6_2341_out0 = v__2831_out1 ? v_MUX5_8840_out0 : v_MUX4_376_out0;
assign v_MUX6_2342_out0 = v__2832_out1 ? v_MUX5_8841_out0 : v_MUX4_377_out0;
assign v_WEN0_2646_out0 = v_WEN0_2588_out0;
assign v_G23_2840_out0 = v_G25_6962_out0 && v_G24_3955_out0;
assign v_G23_2841_out0 = v_G25_6963_out0 && v_G24_3956_out0;
assign v_G2_2891_out0 = v_EXEC1_2634_out0 && v_G3_1720_out0;
assign v_G2_2892_out0 = v_EXEC1_2635_out0 && v_G3_1721_out0;
assign v_G3_2941_out0 = v_FLOAT_7676_out0 && v_NORMAL_13429_out0;
assign v_G3_2942_out0 = v_FLOAT_7677_out0 && v_NORMAL_13430_out0;
assign v_SUB_2957_out0 = v_SUB_8663_out0;
assign v_SUB_2958_out0 = v_SUB_8664_out0;
assign v_G16_3024_out0 = v_EXEC10_8812_out0 && v_REN0_11136_out0;
assign v__3040_out0 = { v__2959_out1,v_BIT_2328_out0 };
assign v_JMI_3212_out0 = v_JMI_13349_out0;
assign v_JMI_3213_out0 = v_JMI_13350_out0;
assign v_CMP_3805_out0 = v_CMP_13609_out0;
assign v_CMP_3806_out0 = v_CMP_13610_out0;
assign v_JEQ_4445_out0 = v_JEQ_2234_out0;
assign v_JEQ_4446_out0 = v_JEQ_2235_out0;
assign v_JUMPADRESS_4745_out0 = v_JUMPADRESS_6964_out0;
assign v_JUMPADRESS_4746_out0 = v_JUMPADRESS_6965_out0;
assign v_SBC_4825_out0 = v_SBC_13605_out0;
assign v_SBC_4826_out0 = v_SBC_13606_out0;
assign v_G2_6884_out0 = v_S_11300_out0 && v_EXEC2_441_out0;
assign v_G2_6885_out0 = v_S_11301_out0 && v_EXEC2_442_out0;
assign v_JMP_7077_out0 = v_JMP_3233_out0;
assign v_JMP_7078_out0 = v_JMP_3234_out0;
assign v_EQ2_7091_out0 = v__4526_out1 == 1'h1;
assign v_EQ2_7092_out0 = v__4527_out1 == 1'h1;
assign v_EXEC2_7181_out0 = v_EXEC2_2647_out0;
assign v_EXEC2_7182_out0 = v_EXEC2_2648_out0;
assign v_TST_8735_out0 = v_TST_3819_out0;
assign v_TST_8736_out0 = v_TST_3820_out0;
assign v_JEQ_8806_out0 = v_JEQ_2234_out0;
assign v_JEQ_8807_out0 = v_JEQ_2235_out0;
assign v_G27_9793_out0 = v__2430_out0 && v_G28_6868_out0;
assign v_G27_9794_out0 = v__2431_out0 && v_G28_6869_out0;
assign v_Wen1_10312_out0 = v_WEN1_8763_out0;
assign v_G7_10332_out0 = v_9_13623_out0 && v_G3_10462_out0;
assign v_G35_10360_out0 = v_STARTBIT_6967_out0 && v_G36_3135_out0;
assign v_G5_10441_out0 = ! v_CMP_13609_out0;
assign v_G5_10442_out0 = ! v_CMP_13610_out0;
assign v_STP_10467_out0 = v_STP_52_out0;
assign v_STP_10468_out0 = v_STP_53_out0;
assign v_MULTI_OPCODE_10797_out0 = v_MULTI_OPCODE_11096_out0;
assign v_MULTI_OPCODE_10798_out0 = v_MULTI_OPCODE_11097_out0;
assign v_UART_10825_out0 = v_UART_1823_out0;
assign v_UART_10826_out0 = v_UART_1824_out0;
assign v__10868_out0 = v__4526_out0[7:0];
assign v__10868_out1 = v__4526_out0[8:1];
assign v__10869_out0 = v__4527_out0[7:0];
assign v__10869_out1 = v__4527_out0[8:1];
assign v_STP_10977_out0 = v_STP_52_out0;
assign v_STP_10978_out0 = v_STP_53_out0;
assign v_G6_11143_out0 = v_G4_1667_out0 && v_NORMAL_181_out0;
assign v_G6_11144_out0 = v_G4_1668_out0 && v_NORMAL_182_out0;
assign v_ADD_11193_out0 = v_ADD_4455_out0;
assign v_ADD_11194_out0 = v_ADD_4456_out0;
assign v_SUB_INSTRUCTION_11195_out0 = v_SUB_INSTRUCTION_2789_out0;
assign v_SUB_INSTRUCTION_11196_out0 = v_SUB_INSTRUCTION_2790_out0;
assign v_BYTERECEIVED_11197_out0 = v_G8_16_out0;
assign v__13253_out0 = v_BIN_5853_out0[3:1];
assign v__13254_out0 = v_BIN_5854_out0[3:1];
assign v_MULTI_INSTRUCTION_13323_out0 = v_MULTI_INSTRUCTION_3953_out0;
assign v_MULTI_INSTRUCTION_13324_out0 = v_MULTI_INSTRUCTION_3954_out0;
assign v_KEXTEND_13329_out0 = v__124_out0;
assign v_KEXTEND_13330_out0 = v__125_out0;
assign v_AND_13556_out0 = v_AND_3858_out0;
assign v_AND_13557_out0 = v_AND_3859_out0;
assign v_ADC_13614_out0 = v_ADC_10393_out0;
assign v_ADC_13615_out0 = v_ADC_10394_out0;
assign v_G3_17_out0 = v_G1_2225_out0 && v_EXEC2_441_out0;
assign v_G3_18_out0 = v_G1_2226_out0 && v_EXEC2_442_out0;
assign v_SR_371_out0 = v_MUX1_534_out0;
assign v_SR_372_out0 = v_MUX1_535_out0;
assign v_TST_409_out0 = v_TST_8735_out0;
assign v_TST_410_out0 = v_TST_8736_out0;
assign v_SR_542_out0 = v_MUX1_534_out0;
assign v_SR_543_out0 = v_MUX1_535_out0;
assign v_MULTI_INSTRUCTION_619_out0 = v_MULTI_INSTRUCTION_13323_out0;
assign v_MULTI_INSTRUCTION_620_out0 = v_MULTI_INSTRUCTION_13324_out0;
assign v_STORE_1195_out0 = v_EQ1_1157_out0;
assign v_STORE_1196_out0 = v_EQ1_1158_out0;
assign v_DOUT1_1207_out0 = v_MUX3_313_out0;
assign v_DOUT1_1208_out0 = v_MUX3_314_out0;
assign v_DOUT2_1733_out0 = v_MUX6_2341_out0;
assign v_DOUT2_1734_out0 = v_MUX6_2342_out0;
assign v_ENABLE_1757_out0 = v_G7_10332_out0;
assign v_STALL_1758_out0 = v_STALL_427_out0;
assign v_STALL_1759_out0 = v_STALL_428_out0;
assign v_ADC_1821_out0 = v_ADC_13614_out0;
assign v_ADC_1822_out0 = v_ADC_13615_out0;
assign v_SR_1956_out0 = v_MUX1_534_out0;
assign v_SR_1957_out0 = v_MUX1_535_out0;
assign v_ENABLE_2018_out0 = v_G35_10360_out0;
assign v_STORE_PCOUNTER_2102_out0 = v_G6_11143_out0;
assign v_STORE_PCOUNTER_2103_out0 = v_G6_11144_out0;
assign v__2146_out0 = { v_C1_10789_out0,v__13253_out0 };
assign v__2147_out0 = { v_C1_10790_out0,v__13254_out0 };
assign v_MUX_ENABLE_2349_out0 = v_G16_3024_out0;
assign v_MULTI_INSTRUCTION_2451_out0 = v_MULTI_INSTRUCTION_13323_out0;
assign v_MULTI_INSTRUCTION_2452_out0 = v_MULTI_INSTRUCTION_13324_out0;
assign v_JMP_2668_out0 = v_JMP_7077_out0;
assign v_JMP_2669_out0 = v_JMP_7078_out0;
assign v_LOAD_3115_out0 = v_EQ2_7091_out0;
assign v_LOAD_3116_out0 = v_EQ2_7092_out0;
assign v_G26_4735_out0 = v_G23_2840_out0 && v__2860_out0;
assign v_G26_4736_out0 = v_G23_2841_out0 && v__2861_out0;
assign v_W_EN_6878_out0 = v__10868_out1;
assign v_W_EN_6879_out0 = v__10869_out1;
assign v_STALL_6910_out0 = v_STALL_427_out0;
assign v_STALL_6911_out0 = v_STALL_428_out0;
assign v__7062_out0 = v__10868_out0[6:0];
assign v__7062_out1 = v__10868_out0[7:1];
assign v__7063_out0 = v__10869_out0[6:0];
assign v__7063_out1 = v__10869_out0[7:1];
assign v_SUB_INSTRUCTION_7085_out0 = v_SUB_INSTRUCTION_11195_out0;
assign v_SUB_INSTRUCTION_7086_out0 = v_SUB_INSTRUCTION_11196_out0;
assign v_WEN1_7716_out0 = v_Wen1_10312_out0;
assign v_CMP_8646_out0 = v_CMP_3805_out0;
assign v_CMP_8647_out0 = v_CMP_3806_out0;
assign v_JMI_8679_out0 = v_JMI_88_out0;
assign v_JMI_8680_out0 = v_JMI_89_out0;
assign v_STP_10307_out0 = v_STP_10977_out0;
assign v_STP_10308_out0 = v_STP_10978_out0;
assign v_AD3_10482_out0 = v_MUX2_1145_out0;
assign v_AD3_10483_out0 = v_MUX2_1146_out0;
assign v_UART_10516_out0 = v_UART_10825_out0;
assign v_UART_10517_out0 = v_UART_10826_out0;
assign v_done_receiving_10604_out0 = v_BYTERECEIVED_11197_out0;
assign v_SR_10607_out0 = v_MUX1_534_out0;
assign v_SR_10608_out0 = v_MUX1_535_out0;
assign v_SBC_11051_out0 = v_SBC_4825_out0;
assign v_SBC_11052_out0 = v_SBC_4826_out0;
assign v_STP_11240_out0 = v_STP_10467_out0;
assign v_STP_11241_out0 = v_STP_10468_out0;
assign v_SUB_12247_out0 = v_SUB_2957_out0;
assign v_SUB_12248_out0 = v_SUB_2958_out0;
assign v_AD3_13272_out0 = v_MUX2_1145_out0;
assign v_AD3_13273_out0 = v_MUX2_1146_out0;
assign v_WEN0_13300_out0 = v_WEN0_2646_out0;
assign v_JEQ_13560_out0 = v_JEQ_4445_out0;
assign v_JEQ_13561_out0 = v_JEQ_4446_out0;
assign v_G1_13776_out0 = v_G2_2891_out0 || v_EXEC2_3241_out0;
assign v_G1_13777_out0 = v_G2_2892_out0 || v_EXEC2_3242_out0;
assign v_LOAD_231_out0 = v_LOAD_3115_out0;
assign v_LOAD_232_out0 = v_LOAD_3116_out0;
assign v_ROR_282_out0 = v_SR_542_out0 == 2'h3;
assign v_ROR_283_out0 = v_SR_543_out0 == 2'h3;
assign v_G6_327_out0 = v_C_3197_out0 && v_ADC_1821_out0;
assign v_G6_328_out0 = v_C_3198_out0 && v_ADC_1822_out0;
assign v_G9_407_out0 = ! v_W_EN_6878_out0;
assign v_G9_408_out0 = ! v_W_EN_6879_out0;
assign v_G9_411_out0 = ((v_AND_13556_out0 && !v_TST_409_out0) || (!v_AND_13556_out0) && v_TST_409_out0);
assign v_G9_412_out0 = ((v_AND_13557_out0 && !v_TST_410_out0) || (!v_AND_13557_out0) && v_TST_410_out0);
assign v_LSR_418_out0 = v_SR_371_out0 == 2'h1;
assign v_LSR_419_out0 = v_SR_372_out0 == 2'h1;
assign v_G5_454_out0 = v_STORE_1195_out0 && v_EXEC1_20_out0;
assign v_G5_455_out0 = v_STORE_1196_out0 && v_EXEC1_21_out0;
assign v_RD_501_out0 = v_DOUT1_1207_out0;
assign v_RD_502_out0 = v_DOUT1_1208_out0;
assign v_STORE_540_out0 = v_STORE_1195_out0;
assign v_STORE_541_out0 = v_STORE_1196_out0;
assign v_ROR_544_out0 = v_SR_371_out0 == 2'h3;
assign v_ROR_545_out0 = v_SR_372_out0 == 2'h3;
assign v_LSR_1174_out0 = v_SR_542_out0 == 2'h1;
assign v_LSR_1175_out0 = v_SR_543_out0 == 2'h1;
assign v_G9_1671_out0 = ! v_STALL_6910_out0;
assign v_G9_1672_out0 = ! v_STALL_6911_out0;
assign v_LSL_1861_out0 = v_SR_542_out0 == 2'h0;
assign v_LSL_1862_out0 = v_SR_543_out0 == 2'h0;
assign v_G2_1887_out0 = v_W_EN_6878_out0 && v_EXEC1_20_out0;
assign v_G2_1888_out0 = v_W_EN_6879_out0 && v_EXEC1_21_out0;
assign v_MUX1_2409_out0 = v_C_379_out0 ? v__2146_out0 : v_BIN_5853_out0;
assign v_MUX1_2410_out0 = v_C_380_out0 ? v__2147_out0 : v_BIN_5854_out0;
assign v_LSL_2842_out0 = v_SR_10607_out0 == 2'h0;
assign v_LSL_2843_out0 = v_SR_10608_out0 == 2'h0;
assign v_STORE_pccounter_2883_out0 = v_STORE_PCOUNTER_2102_out0;
assign v_STORE_pccounter_2884_out0 = v_STORE_PCOUNTER_2103_out0;
assign v_G3_2903_out0 = v_LOAD_3115_out0 && v_EXEC2_7181_out0;
assign v_G3_2904_out0 = v_LOAD_3116_out0 && v_EXEC2_7182_out0;
assign v_G1_3018_out0 = v_SBC_11051_out0 && v_C_3197_out0;
assign v_G1_3019_out0 = v_SBC_11052_out0 && v_C_3198_out0;
assign v_LSL_3047_out0 = v_SR_371_out0 == 2'h0;
assign v_LSL_3048_out0 = v_SR_372_out0 == 2'h0;
assign v_LSL_3182_out0 = v_SR_1956_out0 == 2'h0;
assign v_LSL_3183_out0 = v_SR_1957_out0 == 2'h0;
assign v_ROR_3286_out0 = v_SR_10607_out0 == 2'h3;
assign v_ROR_3287_out0 = v_SR_10608_out0 == 2'h3;
assign v_ROR_3288_out0 = v_SR_1956_out0 == 2'h3;
assign v_ROR_3289_out0 = v_SR_1957_out0 == 2'h3;
assign v_UART_3893_out0 = v_UART_10516_out0;
assign v_UART_3894_out0 = v_UART_10517_out0;
assign v_G5_4477_out0 = v_SUB_12247_out0 || v_CMP_8646_out0;
assign v_G5_4478_out0 = v_SUB_12248_out0 || v_CMP_8647_out0;
assign v_G4_4738_out0 = ((v_SBC_11051_out0 && !v_ADC_1821_out0) || (!v_SBC_11051_out0) && v_ADC_1821_out0);
assign v_G4_4739_out0 = ((v_SBC_11052_out0 && !v_ADC_1822_out0) || (!v_SBC_11052_out0) && v_ADC_1822_out0);
assign v_G29_5834_out0 = v_G26_4735_out0 || v_G27_9793_out0;
assign v_G29_5835_out0 = v_G26_4736_out0 || v_G27_9794_out0;
assign v_LSR_6912_out0 = v_SR_1956_out0 == 2'h1;
assign v_LSR_6913_out0 = v_SR_1957_out0 == 2'h1;
assign v_G3_8665_out0 = ((v_SUB_12247_out0 && !v_CMP_8646_out0) || (!v_SUB_12247_out0) && v_CMP_8646_out0);
assign v_G3_8666_out0 = ((v_SUB_12248_out0 && !v_CMP_8647_out0) || (!v_SUB_12248_out0) && v_CMP_8647_out0);
assign v_AD3_8671_out0 = v_AD3_13272_out0;
assign v_AD3_8672_out0 = v_AD3_13273_out0;
assign v_ASR_8754_out0 = v_SR_1956_out0 == 2'h2;
assign v_ASR_8755_out0 = v_SR_1957_out0 == 2'h2;
assign v_G18_8799_out0 = !(v_ENABLE_2018_out0 || v_Q7_6888_out0);
assign v_STALL_10281_out0 = v_STALL_1758_out0;
assign v_STALL_10282_out0 = v_STALL_1759_out0;
assign v_G4_10283_out0 = v_G5_10914_out0 && v_STALL_6910_out0;
assign v_G4_10284_out0 = v_G5_10915_out0 && v_STALL_6911_out0;
assign v_G19_10327_out0 = ! v_STP_11240_out0;
assign v_G19_10328_out0 = ! v_STP_11241_out0;
assign v_ASR_10366_out0 = v_SR_542_out0 == 2'h2;
assign v_ASR_10367_out0 = v_SR_543_out0 == 2'h2;
assign v_RX_DONE_RECEIVING_10484_out0 = v_done_receiving_10604_out0;
assign v__10490_out0 = v__7062_out0[5:0];
assign v__10490_out1 = v__7062_out0[6:1];
assign v__10491_out0 = v__7063_out0[5:0];
assign v__10491_out1 = v__7063_out0[6:1];
assign v_ASR_10566_out0 = v_SR_371_out0 == 2'h2;
assign v_ASR_10567_out0 = v_SR_372_out0 == 2'h2;
assign v_P_10682_out0 = v__7062_out1;
assign v_P_10683_out0 = v__7063_out1;
assign v_G17_10710_out0 = v_MUX_ENABLE_2349_out0 && v_G18_567_out0;
assign v_WENMULTI_11206_out0 = v_G1_13776_out0;
assign v_WENMULTI_11207_out0 = v_G1_13777_out0;
assign v_G4_12243_out0 = v_G5_10441_out0 && v_G3_17_out0;
assign v_G4_12244_out0 = v_G5_10442_out0 && v_G3_18_out0;
assign v_MULTI_INSTRUCTION_13308_out0 = v_MULTI_INSTRUCTION_619_out0;
assign v_MULTI_INSTRUCTION_13309_out0 = v_MULTI_INSTRUCTION_620_out0;
assign v_LSR_13331_out0 = v_SR_10607_out0 == 2'h1;
assign v_LSR_13332_out0 = v_SR_10608_out0 == 2'h1;
assign v_G11_13439_out0 = v_G20_598_out0 || v_STP_11240_out0;
assign v_G11_13440_out0 = v_G20_599_out0 || v_STP_11241_out0;
assign v_RM_13597_out0 = v_DOUT2_1733_out0;
assign v_RM_13598_out0 = v_DOUT2_1734_out0;
assign v_ASR_13713_out0 = v_SR_10607_out0 == 2'h2;
assign v_ASR_13714_out0 = v_SR_10608_out0 == 2'h2;
assign v_RM_13750_out0 = v_DOUT2_1733_out0;
assign v_RM_13751_out0 = v_DOUT2_1734_out0;
assign v_G30_184_out0 = v_G2_1888_out0 && v_STALL_DUAL_CORE_12235_out0;
assign v__1140_out0 = v__10490_out0[1:0];
assign v__1140_out1 = v__10490_out0[5:4];
assign v__1141_out0 = v__10491_out0[1:0];
assign v__1141_out1 = v__10491_out0[5:4];
assign v_G1_1191_out0 = ! v__10490_out1;
assign v_G1_1192_out0 = ! v__10491_out1;
assign v_G8_1765_out0 = v_G7_1684_out0 || v_G4_10283_out0;
assign v_G8_1766_out0 = v_G7_1685_out0 || v_G4_10284_out0;
assign v_G22_1900_out0 = v_G11_13440_out0 && v_STALL_DUAL_CORE_4696_out0;
assign v_WEN_MULTI_2388_out0 = v_WENMULTI_11206_out0;
assign v_WEN_MULTI_2389_out0 = v_WENMULTI_11207_out0;
assign v_G11_2626_out0 = v_G5_10914_out0 && v_G9_1671_out0;
assign v_G11_2627_out0 = v_G5_10915_out0 && v_G9_1672_out0;
assign v_RDOUT_2787_out0 = v_RD_501_out0;
assign v_RDOUT_2788_out0 = v_RD_502_out0;
assign v_LOAD_2899_out0 = v_LOAD_231_out0;
assign v_LOAD_2900_out0 = v_LOAD_232_out0;
assign v_DONE_RECEIVING_3084_out0 = v_RX_DONE_RECEIVING_10484_out0;
assign v_RXBYTERECEIVED_3269_out0 = v_RX_DONE_RECEIVING_10484_out0;
assign v_G21_3808_out0 = v_G18_8799_out0 || v_G22_10983_out0;
assign v_RD_3891_out0 = v_RD_501_out0;
assign v_RD_3892_out0 = v_RD_502_out0;
assign v_OP1_3899_out0 = v_RD_501_out0;
assign v_OP1_3900_out0 = v_RD_502_out0;
assign v_G8_4453_out0 = v_G1_3018_out0 || v_G6_327_out0;
assign v_G8_4454_out0 = v_G1_3019_out0 || v_G6_328_out0;
assign v_G7_4474_out0 = v_P_10682_out0 && v_EXEC1_20_out0;
assign v_G7_4475_out0 = v_P_10683_out0 && v_EXEC1_21_out0;
assign v_G10_4479_out0 = v_EXEC2_7181_out0 && v_P_10682_out0;
assign v_G10_4480_out0 = v_EXEC2_7182_out0 && v_P_10683_out0;
assign v_RM_4537_out0 = v_RM_13750_out0;
assign v_RM_4538_out0 = v_RM_13751_out0;
assign v_STORE_WEN_4544_out0 = v_STORE_pccounter_2883_out0;
assign v_STORE_WEN_4545_out0 = v_STORE_pccounter_2884_out0;
assign v_EN_4593_out0 = v_G29_5834_out0;
assign v_EN_4594_out0 = v_G29_5835_out0;
assign v_G24_4780_out0 = ! v_G17_10710_out0;
assign v_G5_7106_out0 = v_MULTI_INSTRUCTION_13308_out0 || v_DIV_INSTRUCTION_4614_out0;
assign v_G5_7107_out0 = v_MULTI_INSTRUCTION_13309_out0 || v_DIV_INSTRUCTION_4615_out0;
assign v_RM_8731_out0 = v_RM_13750_out0;
assign v_RM_8732_out0 = v_RM_13751_out0;
assign v_MUX1_8813_out0 = v_C_8653_out0 ? v_KEXTEND_13329_out0 : v_RM_13597_out0;
assign v_MUX1_8814_out0 = v_C_8654_out0 ? v_KEXTEND_13330_out0 : v_RM_13598_out0;
assign v_MUX10_10395_out0 = v_MULTI_INSTRUCTION_13308_out0 ? v_C13_405_out0 : v_C12_2113_out0;
assign v_MUX10_10396_out0 = v_MULTI_INSTRUCTION_13309_out0 ? v_C13_406_out0 : v_C12_2114_out0;
assign v_RAMWEN_10701_out0 = v_G5_454_out0;
assign v_RAMWEN_10702_out0 = v_G5_455_out0;
assign v_B_10793_out0 = v_MUX1_2409_out0;
assign v_B_10794_out0 = v_MUX1_2410_out0;
assign v_STORE_10831_out0 = v_STORE_540_out0;
assign v_STORE_10832_out0 = v_STORE_541_out0;
assign v_WENALU_10866_out0 = v_G4_12243_out0;
assign v_WENALU_10867_out0 = v_G4_12244_out0;
assign v_UART_11128_out0 = v_UART_3893_out0;
assign v_UART_11129_out0 = v_UART_3894_out0;
assign v_G2_11134_out0 = ((v_ADD_11193_out0 && !v_G3_8665_out0) || (!v_ADD_11193_out0) && v_G3_8665_out0);
assign v_G2_11135_out0 = ((v_ADD_11194_out0 && !v_G3_8666_out0) || (!v_ADD_11194_out0) && v_G3_8666_out0);
assign v_G11_11165_out0 = v_G5_4477_out0 || v_SBC_11051_out0;
assign v_G11_11166_out0 = v_G5_4478_out0 || v_SBC_11052_out0;
assign v_RM_11167_out0 = v_RM_13750_out0;
assign v_RM_11168_out0 = v_RM_13751_out0;
assign v_G4_13702_out0 = ! v_MULTI_INSTRUCTION_13308_out0;
assign v_G4_13703_out0 = ! v_MULTI_INSTRUCTION_13309_out0;
assign v_EN_STALL_13747_out0 = v_G17_10710_out0;
assign v_RXBYTERECEIVED_91_out0 = v_RXBYTERECEIVED_3269_out0;
assign v_SEL6_103_out0 = v_RM_11167_out0[9:0];
assign v_SEL6_104_out0 = v_RM_11168_out0[9:0];
assign v_G10_130_out0 = v_G8_4453_out0 || v_G5_4477_out0;
assign v_G10_131_out0 = v_G8_4454_out0 || v_G5_4478_out0;
assign v_G7_169_out0 = ((v_G2_11134_out0 && !v_G4_4738_out0) || (!v_G2_11134_out0) && v_G4_4738_out0);
assign v_G7_170_out0 = ((v_G2_11135_out0 && !v_G4_4739_out0) || (!v_G2_11135_out0) && v_G4_4739_out0);
assign v__186_out0 = v_B_10793_out0[3:3];
assign v__187_out0 = v_B_10794_out0[3:3];
assign v_G4_220_out0 = v_G30_184_out0 || v_G3_2904_out0;
assign v__413_out0 = v_B_10793_out0[1:1];
assign v__414_out0 = v_B_10794_out0[1:1];
assign v__1728_out0 = v_B_10793_out0[0:0];
assign v__1729_out0 = v_B_10794_out0[0:0];
assign v_WENRAM_2326_out0 = v_RAMWEN_10701_out0;
assign v_WENRAM_2327_out0 = v_RAMWEN_10702_out0;
assign v_G18_2407_out0 = v_G16_2310_out0 && v_G8_1765_out0;
assign v_G18_2408_out0 = v_G16_2311_out0 && v_G8_1766_out0;
assign v_RM_2432_out0 = v_RM_8731_out0;
assign v_RM_2433_out0 = v_RM_8732_out0;
assign v_SEL3_2615_out0 = v_RD_3891_out0[15:15];
assign v_SEL3_2616_out0 = v_RD_3892_out0[15:15];
assign v_G8_2623_out0 = v_G9_407_out0 && v_G10_4479_out0;
assign v_G8_2624_out0 = v_G9_408_out0 && v_G10_4480_out0;
assign v_SUB_2910_out0 = v_G22_1900_out0;
assign v_SEL1_2917_out0 = v_RD_3891_out0[14:10];
assign v_SEL1_2918_out0 = v_RD_3892_out0[14:10];
assign v_OP1_2979_out0 = v_OP1_3899_out0;
assign v_OP1_2980_out0 = v_OP1_3900_out0;
assign v_G23_3083_out0 = v_WEN1_7716_out0 && v_G24_4780_out0;
assign v_SUB_4616_out0 = v_G11_11165_out0;
assign v_SUB_4618_out0 = v_G11_11166_out0;
assign v_M_4701_out0 = v__1140_out0;
assign v_M_4702_out0 = v__1141_out0;
assign v_DONE_RECEIVING_5857_out0 = v_DONE_RECEIVING_3084_out0;
assign v_LOAD_7110_out0 = v_LOAD_2899_out0;
assign v_LOAD_7111_out0 = v_LOAD_2900_out0;
assign v_SEL4_7636_out0 = v_RM_11167_out0[15:15];
assign v_SEL4_7637_out0 = v_RM_11168_out0[15:15];
assign v_N_7642_out0 = v__1140_out1;
assign v_N_7643_out0 = v__1141_out1;
assign v_WENALU_8659_out0 = v_WENALU_10866_out0;
assign v_WENALU_8660_out0 = v_WENALU_10867_out0;
assign v_SEL5_8767_out0 = v_RD_3891_out0[9:0];
assign v_SEL5_8768_out0 = v_RD_3892_out0[9:0];
assign v_REGISTER_OUT_10268_out0 = v_RDOUT_2787_out0;
assign v_REGISTER_OUT_10269_out0 = v_RDOUT_2788_out0;
assign v_G12_10321_out0 = v_G11_2626_out0 && v_G2_6791_out0;
assign v_G12_10322_out0 = v_G11_2627_out0 && v_G2_6792_out0;
assign v_EN_STALL_10344_out0 = v_EN_STALL_13747_out0;
assign v_WEN_MULTI_10381_out0 = v_WEN_MULTI_2388_out0;
assign v_WEN_MULTI_10382_out0 = v_WEN_MULTI_2389_out0;
assign v_U_10469_out0 = v_G1_1191_out0;
assign v_U_10470_out0 = v_G1_1192_out0;
assign v__10785_out0 = v_B_10793_out0[2:2];
assign v__10786_out0 = v_B_10794_out0[2:2];
assign v_IN_11258_out0 = v_MUX1_8813_out0;
assign v_IN_11259_out0 = v_MUX1_8814_out0;
assign v_STORE_13298_out0 = v_STORE_10831_out0;
assign v_STORE_13299_out0 = v_STORE_10832_out0;
assign v_SEL2_13327_out0 = v_RM_11167_out0[14:10];
assign v_SEL2_13328_out0 = v_RM_11168_out0[14:10];
assign v_RM_13508_out0 = v_RM_4537_out0;
assign v_RM_13509_out0 = v_RM_4538_out0;
assign v_WEN_MULTI_35_out0 = v_WEN_MULTI_10381_out0;
assign v_WEN_MULTI_36_out0 = v_WEN_MULTI_10382_out0;
assign v_IN_98_out0 = v_IN_11258_out0;
assign v_IN_99_out0 = v_IN_11259_out0;
assign v_STORE_221_out0 = v_STORE_13298_out0;
assign v_STORE_222_out0 = v_STORE_13299_out0;
assign v_G5_230_out0 = ((v__3271_out0 && !v_SUB_2910_out0) || (!v__3271_out0) && v_SUB_2910_out0);
assign v_RAM_IN_233_out0 = v_REGISTER_OUT_10268_out0;
assign v_RAM_IN_234_out0 = v_REGISTER_OUT_10269_out0;
assign v_RD_SIGN_285_out0 = v_SEL3_2615_out0;
assign v_RD_SIGN_286_out0 = v_SEL3_2616_out0;
assign v_G10_1755_out0 = v_G6_2905_out0 || v_G12_10321_out0;
assign v_G10_1756_out0 = v_G6_2906_out0 || v_G12_10322_out0;
assign v_RD_SIG_1769_out0 = v_SEL5_8767_out0;
assign v_RD_SIG_1770_out0 = v_SEL5_8768_out0;
assign v_G17_1903_out0 = v_RXBYTERECEIVED_91_out0 && v_Q1_3993_out0;
assign v_G8_2025_out0 = ((v__172_out0 && !v_SUB_2910_out0) || (!v__172_out0) && v_SUB_2910_out0);
assign v_OP1_2060_out0 = v_OP1_2979_out0;
assign v_OP1_2061_out0 = v_OP1_2980_out0;
assign v_EN_2330_out0 = v__1728_out0;
assign v_EN_2331_out0 = v__1729_out0;
assign v_G9_2333_out0 = ((v__2269_out0 && !v_SUB_2910_out0) || (!v__2269_out0) && v_SUB_2910_out0);
assign v_G6_2417_out0 = ((v__2023_out0 && !v_SUB_2910_out0) || (!v__2023_out0) && v_SUB_2910_out0);
assign v_EN_2445_out0 = v__186_out0;
assign v_EN_2446_out0 = v__187_out0;
assign v_OP2_EXP_2548_out0 = v_SEL2_13327_out0;
assign v_OP2_EXP_2549_out0 = v_SEL2_13328_out0;
assign v_G11_2551_out0 = ((v__61_out0 && !v_SUB_2910_out0) || (!v__61_out0) && v_SUB_2910_out0);
assign v_G3_2622_out0 = ((v__288_out0 && !v_SUB_2910_out0) || (!v__288_out0) && v_SUB_2910_out0);
assign v_G10_2633_out0 = ((v__11243_out0 && !v_SUB_2910_out0) || (!v__11243_out0) && v_SUB_2910_out0);
assign v__3035_out0 = v_RM_13508_out0[11:0];
assign v__3035_out1 = v_RM_13508_out0[15:4];
assign v__3036_out0 = v_RM_13509_out0[11:0];
assign v__3036_out1 = v_RM_13509_out0[15:4];
assign v_G2_3240_out0 = ((v__3124_out0 && !v_SUB_2910_out0) || (!v__3124_out0) && v_SUB_2910_out0);
assign v_G19_3860_out0 = v_RXBYTERECEIVED_91_out0 || v_Q1_3993_out0;
assign v_SUB_4617_out0 = v_U_10469_out0;
assign v_SUB_4619_out0 = v_U_10470_out0;
assign v_WENRAM_4650_out0 = v_WENRAM_2326_out0;
assign v_WENRAM_4651_out0 = v_WENRAM_2327_out0;
assign v_G12_4700_out0 = ((v__1876_out0 && !v_SUB_2910_out0) || (!v__1876_out0) && v_SUB_2910_out0);
assign v_G7_4822_out0 = ((v__13397_out0 && !v_SUB_2910_out0) || (!v__13397_out0) && v_SUB_2910_out0);
assign v_byte_ready_5843_out0 = v_DONE_RECEIVING_5857_out0;
assign v_LOAD_8765_out0 = v_LOAD_7110_out0;
assign v_LOAD_8766_out0 = v_LOAD_7111_out0;
assign v_RD_EXP_8846_out0 = v_SEL1_2917_out0;
assign v_RD_EXP_8847_out0 = v_SEL1_2918_out0;
assign v_EN_10474_out0 = v__413_out0;
assign v_EN_10475_out0 = v__414_out0;
assign v_G1_10478_out0 = ((v__13563_out0 && !v_SUB_2910_out0) || (!v__13563_out0) && v_SUB_2910_out0);
assign v_G21_10788_out0 = v_G23_3083_out0 || v_WEN0_13300_out0;
assign v_OP2_SIGN_10839_out0 = v_SEL4_7636_out0;
assign v_OP2_SIGN_10840_out0 = v_SEL4_7637_out0;
assign v__11229_out0 = { v_N_7642_out0,v_C1_3210_out0 };
assign v__11230_out0 = { v_N_7643_out0,v_C1_3211_out0 };
assign v_G4_12239_out0 = ((v__180_out0 && !v_SUB_2910_out0) || (!v__180_out0) && v_SUB_2910_out0);
assign v_EN_13181_out0 = v__10785_out0;
assign v_EN_13182_out0 = v__10786_out0;
assign v_G6_13258_out0 = v_G8_2623_out0 || v_G7_4474_out0;
assign v_G6_13259_out0 = v_G8_2624_out0 || v_G7_4475_out0;
assign v_OP2_SIG_13301_out0 = v_SEL6_103_out0;
assign v_OP2_SIG_13302_out0 = v_SEL6_104_out0;
assign v_STALL_DUAL_CORE_13617_out0 = v_EN_STALL_10344_out0;
assign v_WENLDST_13756_out0 = v_G4_220_out0;
assign v_OP2_EXP_536_out0 = v_OP2_EXP_2548_out0;
assign v_OP2_EXP_537_out0 = v_OP2_EXP_2549_out0;
assign v__1708_out0 = { v_G1_10478_out0,v_G2_3240_out0 };
assign v_SIG_RM_1767_out0 = v_OP2_SIG_13301_out0;
assign v_SIG_RM_1768_out0 = v_OP2_SIG_13302_out0;
assign v_RD_SIGN_2405_out0 = v_RD_SIGN_285_out0;
assign v_RD_SIGN_2406_out0 = v_RD_SIGN_286_out0;
assign v_WENLDST_2683_out0 = v_WENLDST_13756_out0;
assign v_WEN_3204_out0 = v_G21_10788_out0;
assign v_LOAD_3949_out0 = v_LOAD_8765_out0;
assign v_LOAD_3950_out0 = v_LOAD_8766_out0;
assign v_RD_EXP_3951_out0 = v_RD_EXP_8846_out0;
assign v_RD_EXP_3952_out0 = v_RD_EXP_8847_out0;
assign v_G2_4467_out0 = ! v_STALL_DUAL_CORE_13617_out0;
assign v_EXP_RM_4743_out0 = v_OP2_EXP_2548_out0;
assign v_EXP_RM_4744_out0 = v_OP2_EXP_2549_out0;
assign v__4831_out0 = v_IN_98_out0[14:0];
assign v__4831_out1 = v_IN_98_out0[15:1];
assign v__4832_out0 = v_IN_99_out0[14:0];
assign v__4832_out1 = v_IN_99_out0[15:1];
assign v_EXP_RD_5855_out0 = v_RD_EXP_8846_out0;
assign v_EXP_RD_5856_out0 = v_RD_EXP_8847_out0;
assign v_A_10275_out0 = v_OP1_2060_out0;
assign v_A_10277_out0 = v_OP1_2061_out0;
assign v_BYTE_READY_11173_out0 = v_byte_ready_5843_out0;
assign v_OP2_SIGN_11208_out0 = v_OP2_SIGN_10839_out0;
assign v_OP2_SIGN_11209_out0 = v_OP2_SIGN_10840_out0;
assign v_A_11251_out0 = v__11229_out0;
assign v_A_11253_out0 = v__11230_out0;
assign v_SIG_RD_11298_out0 = v_RD_SIG_1769_out0;
assign v_SIG_RD_11299_out0 = v_RD_SIG_1770_out0;
assign v_G14_13268_out0 = v_G10_1755_out0 || v_G13_7083_out0;
assign v_G14_13269_out0 = v_G10_1756_out0 || v_G13_7084_out0;
assign v_UNUSED_13431_out0 = v__3035_out1;
assign v_UNUSED_13432_out0 = v__3036_out1;
assign v_IN_13788_out0 = v_IN_98_out0;
assign v_IN_13789_out0 = v_IN_99_out0;
assign v__1_out0 = v_A_10275_out0[4:4];
assign v__3_out0 = v_A_10277_out0[4:4];
assign v__78_out0 = v_A_11251_out0[3:3];
assign v__80_out0 = v_A_11253_out0[3:3];
assign v__193_out0 = v_A_11251_out0[15:15];
assign v__195_out0 = v_A_11253_out0[15:15];
assign v_G1_289_out0 = ((v_OP2_SIGN_11208_out0 && !v_SUB_INSTRUCTION_7085_out0) || (!v_OP2_SIGN_11208_out0) && v_SUB_INSTRUCTION_7085_out0);
assign v_G1_290_out0 = ((v_OP2_SIGN_11209_out0 && !v_SUB_INSTRUCTION_7086_out0) || (!v_OP2_SIGN_11209_out0) && v_SUB_INSTRUCTION_7086_out0);
assign v__322_out0 = v_A_11251_out0[0:0];
assign v__324_out0 = v_A_11253_out0[0:0];
assign v__330_out0 = v_A_11251_out0[9:9];
assign v__332_out0 = v_A_11253_out0[9:9];
assign v_WENLS_601_out0 = v_WENLDST_2683_out0;
assign v__1693_out0 = v_A_10275_out0[5:5];
assign v__1695_out0 = v_A_10277_out0[5:5];
assign v__1748_out0 = v_A_10275_out0[11:11];
assign v__1750_out0 = v_A_10277_out0[11:11];
assign v__1894_out0 = v_A_10275_out0[0:0];
assign v__1896_out0 = v_A_10277_out0[0:0];
assign v__2094_out0 = v_A_11251_out0[13:13];
assign v__2096_out0 = v_A_11253_out0[13:13];
assign v__2151_out0 = v_A_10275_out0[2:2];
assign v__2153_out0 = v_A_10277_out0[2:2];
assign v_WEN_2154_out0 = v_WEN_3204_out0;
assign v__2387_out0 = { v__1708_out0,v_G3_2622_out0 };
assign v__2419_out0 = v_A_11251_out0[6:6];
assign v__2421_out0 = v_A_11253_out0[6:6];
assign v_RD_EXP_2601_out0 = v_RD_EXP_3951_out0;
assign v_RD_EXP_2602_out0 = v_RD_EXP_3952_out0;
assign v__2761_out0 = v_A_10275_out0[15:15];
assign v__2763_out0 = v_A_10277_out0[15:15];
assign v__2876_out0 = v_A_10275_out0[12:12];
assign v__2878_out0 = v_A_10277_out0[12:12];
assign v__2880_out0 = v_A_10275_out0[3:3];
assign v__2882_out0 = v_A_10277_out0[3:3];
assign v__3120_out0 = v_A_11251_out0[14:14];
assign v__3122_out0 = v_A_11253_out0[14:14];
assign v_STALL_DUAL_CORE_3127_out0 = v_G2_4467_out0;
assign v__3248_out0 = v_A_10275_out0[8:8];
assign v__3250_out0 = v_A_10277_out0[8:8];
assign v__3283_out0 = v_A_11251_out0[2:2];
assign v__3285_out0 = v_A_11253_out0[2:2];
assign v__4598_out0 = v_A_10275_out0[10:10];
assign v__4600_out0 = v_A_10277_out0[10:10];
assign v__4712_out0 = v_A_10275_out0[13:13];
assign v__4714_out0 = v_A_10277_out0[13:13];
assign v_BYTE_READY_7022_out0 = v_BYTE_READY_11173_out0;
assign v__7179_out0 = { v_C1_604_out0,v__4831_out0 };
assign v__7180_out0 = { v_C1_605_out0,v__4832_out0 };
assign v__8749_out0 = v_A_11251_out0[8:8];
assign v__8751_out0 = v_A_11253_out0[8:8];
assign v_MUX3_8818_out0 = v_IR15_2465_out0 ? v_WENALU_8660_out0 : v_WENLDST_2683_out0;
assign v__8828_out0 = v_A_11251_out0[7:7];
assign v__8830_out0 = v_A_11253_out0[7:7];
assign v__8849_out0 = v_A_10275_out0[14:14];
assign v__8851_out0 = v_A_10277_out0[14:14];
assign v_EQ2_10347_out0 = v_EXP_RM_4743_out0 == 5'h0;
assign v_EQ2_10348_out0 = v_EXP_RM_4744_out0 == 5'h0;
assign v__10378_out0 = v_A_11251_out0[5:5];
assign v__10380_out0 = v_A_11253_out0[5:5];
assign v_OP2_EXP_10383_out0 = v_OP2_EXP_536_out0;
assign v_OP2_EXP_10384_out0 = v_OP2_EXP_537_out0;
assign v__10386_out0 = v_A_11251_out0[1:1];
assign v__10388_out0 = v_A_11253_out0[1:1];
assign v__10696_out0 = v_A_11251_out0[4:4];
assign v__10698_out0 = v_A_11253_out0[4:4];
assign v__10778_out0 = v_A_11251_out0[12:12];
assign v__10780_out0 = v_A_11253_out0[12:12];
assign v__10863_out0 = v_A_11251_out0[10:10];
assign v__10865_out0 = v_A_11253_out0[10:10];
assign v__11057_out0 = { v_G14_13268_out0,v_G18_2407_out0 };
assign v__11058_out0 = { v_G14_13269_out0,v_G18_2408_out0 };
assign v__11150_out0 = v_A_10275_out0[6:6];
assign v__11152_out0 = v_A_10277_out0[6:6];
assign v_UNNOTUSED_11220_out0 = v__4831_out1;
assign v_UNNOTUSED_11221_out0 = v__4832_out1;
assign v__13385_out0 = v_A_10275_out0[7:7];
assign v__13387_out0 = v_A_10277_out0[7:7];
assign v_EQ1_13433_out0 = v_EXP_RD_5855_out0 == 5'h0;
assign v_EQ1_13434_out0 = v_EXP_RD_5856_out0 == 5'h0;
assign v__13513_out0 = v_A_10275_out0[1:1];
assign v__13515_out0 = v_A_10277_out0[1:1];
assign v__13553_out0 = v_A_11251_out0[11:11];
assign v__13555_out0 = v_A_11253_out0[11:11];
assign v__13628_out0 = v_A_10275_out0[9:9];
assign v__13630_out0 = v_A_10277_out0[9:9];
assign v_MUX1_31_out0 = v_LSL_3182_out0 ? v__7179_out0 : v_IN_13788_out0;
assign v_MUX1_32_out0 = v_LSL_3183_out0 ? v__7180_out0 : v_IN_13789_out0;
assign v_G3_207_out0 = ((v__3283_out0 && !v_SUB_4617_out0) || (!v__3283_out0) && v_SUB_4617_out0);
assign v_G3_209_out0 = ((v__3285_out0 && !v_SUB_4619_out0) || (!v__3285_out0) && v_SUB_4619_out0);
assign v_D_623_out0 = v__11057_out0;
assign v_D_624_out0 = v__11058_out0;
assign v_G1_646_out0 = ! v_EQ1_13433_out0;
assign v_G1_647_out0 = ! v_EQ1_13434_out0;
assign v_G8_1216_out0 = ((v__8828_out0 && !v_SUB_4617_out0) || (!v__8828_out0) && v_SUB_4617_out0);
assign v_G8_1218_out0 = ((v__8830_out0 && !v_SUB_4619_out0) || (!v__8830_out0) && v_SUB_4619_out0);
assign v_STALL_DUAL_CORE_1738_out0 = v_STALL_DUAL_CORE_3127_out0;
assign v_EQ2_1753_out0 = v_OP2_EXP_10383_out0 == 5'h0;
assign v_EQ2_1754_out0 = v_OP2_EXP_10384_out0 == 5'h0;
assign v_G15_1815_out0 = ((v__3120_out0 && !v_SUB_4617_out0) || (!v__3120_out0) && v_SUB_4617_out0);
assign v_G15_1817_out0 = ((v__3122_out0 && !v_SUB_4619_out0) || (!v__3122_out0) && v_SUB_4619_out0);
assign v_EQ1_2597_out0 = v_RD_EXP_2601_out0 == 5'h0;
assign v_EQ1_2598_out0 = v_RD_EXP_2602_out0 == 5'h0;
assign v_G7_2780_out0 = ((v__2419_out0 && !v_SUB_4617_out0) || (!v__2419_out0) && v_SUB_4617_out0);
assign v_G7_2782_out0 = ((v__2421_out0 && !v_SUB_4619_out0) || (!v__2421_out0) && v_SUB_4619_out0);
assign v__2969_out0 = { v__2387_out0,v_G4_12239_out0 };
assign v_STALL_DUAL_CORE_3264_out0 = v_STALL_DUAL_CORE_3127_out0;
assign v_G12_3346_out0 = ((v__13553_out0 && !v_SUB_4617_out0) || (!v__13553_out0) && v_SUB_4617_out0);
assign v_G12_3348_out0 = ((v__13555_out0 && !v_SUB_4619_out0) || (!v__13555_out0) && v_SUB_4619_out0);
assign v_G14_4534_out0 = ((v__2094_out0 && !v_SUB_4617_out0) || (!v__2094_out0) && v_SUB_4617_out0);
assign v_G14_4536_out0 = ((v__2096_out0 && !v_SUB_4619_out0) || (!v__2096_out0) && v_SUB_4619_out0);
assign v_G13_4706_out0 = ((v__10778_out0 && !v_SUB_4617_out0) || (!v__10778_out0) && v_SUB_4617_out0);
assign v_G13_4708_out0 = ((v__10780_out0 && !v_SUB_4619_out0) || (!v__10780_out0) && v_SUB_4619_out0);
assign v_G2_7015_out0 = ! v_EQ2_10347_out0;
assign v_G2_7016_out0 = ! v_EQ2_10348_out0;
assign v_G2_7026_out0 = ((v__10386_out0 && !v_SUB_4617_out0) || (!v__10386_out0) && v_SUB_4617_out0);
assign v_G2_7028_out0 = ((v__10388_out0 && !v_SUB_4619_out0) || (!v__10388_out0) && v_SUB_4619_out0);
assign v_MUX6_8758_out0 = v_MULTI_OPCODE_3021_out0 ? v_WEN_MULTI_2389_out0 : v_MUX3_8818_out0;
assign v_BYTE_READY_10559_out0 = v_BYTE_READY_7022_out0;
assign v_G5_10569_out0 = ((v__10696_out0 && !v_SUB_4617_out0) || (!v__10696_out0) && v_SUB_4617_out0);
assign v_G5_10571_out0 = ((v__10698_out0 && !v_SUB_4619_out0) || (!v__10698_out0) && v_SUB_4619_out0);
assign v_G4_10998_out0 = ((v__78_out0 && !v_SUB_4617_out0) || (!v__78_out0) && v_SUB_4617_out0);
assign v_G4_11000_out0 = ((v__80_out0 && !v_SUB_4619_out0) || (!v__80_out0) && v_SUB_4619_out0);
assign v_G16_11035_out0 = ((v__193_out0 && !v_SUB_4617_out0) || (!v__193_out0) && v_SUB_4617_out0);
assign v_G16_11037_out0 = ((v__195_out0 && !v_SUB_4619_out0) || (!v__195_out0) && v_SUB_4619_out0);
assign v_WENLS_11261_out0 = v_WENLS_601_out0;
assign v_G10_13216_out0 = ((v__330_out0 && !v_SUB_4617_out0) || (!v__330_out0) && v_SUB_4617_out0);
assign v_G10_13218_out0 = ((v__332_out0 && !v_SUB_4619_out0) || (!v__332_out0) && v_SUB_4619_out0);
assign v_G9_13286_out0 = ((v__8749_out0 && !v_SUB_4617_out0) || (!v__8749_out0) && v_SUB_4617_out0);
assign v_G9_13288_out0 = ((v__8751_out0 && !v_SUB_4619_out0) || (!v__8751_out0) && v_SUB_4619_out0);
assign v_G11_13343_out0 = ((v__10863_out0 && !v_SUB_4617_out0) || (!v__10863_out0) && v_SUB_4617_out0);
assign v_G11_13345_out0 = ((v__10865_out0 && !v_SUB_4619_out0) || (!v__10865_out0) && v_SUB_4619_out0);
assign v_G6_13638_out0 = ((v__10378_out0 && !v_SUB_4617_out0) || (!v__10378_out0) && v_SUB_4617_out0);
assign v_G6_13640_out0 = ((v__10380_out0 && !v_SUB_4619_out0) || (!v__10380_out0) && v_SUB_4619_out0);
assign v_G1_13758_out0 = ((v__322_out0 && !v_SUB_4617_out0) || (!v__322_out0) && v_SUB_4617_out0);
assign v_G1_13760_out0 = ((v__324_out0 && !v_SUB_4619_out0) || (!v__324_out0) && v_SUB_4619_out0);
assign v_WWNELS0_385_out0 = v_WENLS_11261_out0;
assign v_WEN3_1691_out0 = v_MUX6_8758_out0;
assign v__1952_out0 = { v_G1_13758_out0,v_G2_7026_out0 };
assign v__1954_out0 = { v_G1_13760_out0,v_G2_7028_out0 };
assign v_STALL_DUAL_CORE_1958_out0 = v_STALL_DUAL_CORE_1738_out0;
assign v__2771_out0 = { v_SIG_RM_1767_out0,v_G2_7015_out0 };
assign v__2772_out0 = { v_SIG_RM_1768_out0,v_G2_7016_out0 };
assign v_BYTE_READY_2853_out0 = v_BYTE_READY_10559_out0;
assign v__4605_out0 = v_D_623_out0[0:0];
assign v__4605_out1 = v_D_623_out0[1:1];
assign v__4606_out0 = v_D_624_out0[0:0];
assign v__4606_out1 = v_D_624_out0[1:1];
assign v_STALL_DUAL_CORE_4695_out0 = v_STALL_DUAL_CORE_1738_out0;
assign v__4856_out0 = v_MUX1_31_out0[0:0];
assign v__4856_out1 = v_MUX1_31_out0[15:15];
assign v__4857_out0 = v_MUX1_32_out0[0:0];
assign v__4857_out1 = v_MUX1_32_out0[15:15];
assign v__5850_out0 = { v__2969_out0,v_G5_230_out0 };
assign v__7714_out0 = { v_SIG_RD_11298_out0,v_G1_646_out0 };
assign v__7715_out0 = { v_SIG_RD_11299_out0,v_G1_647_out0 };
assign v_STALL_DUAL_CORE_12234_out0 = v_STALL_DUAL_CORE_3264_out0;
assign v_MUX13_13647_out0 = v_EQ1_2597_out0 ? v_0B00001_10554_out0 : v_RD_EXP_2601_out0;
assign v_MUX13_13648_out0 = v_EQ1_2598_out0 ? v_0B00001_10555_out0 : v_RD_EXP_2602_out0;
assign v_MUX12_13783_out0 = v_EQ2_1753_out0 ? v_0B00001_10554_out0 : v_OP2_EXP_10383_out0;
assign v_MUX12_13784_out0 = v_EQ2_1754_out0 ? v_0B00001_10555_out0 : v_OP2_EXP_10384_out0;
assign v__97_out0 = { v__5850_out0,v_G6_2417_out0 };
assign v_G30_183_out0 = v_G2_1887_out0 && v_STALL_DUAL_CORE_12234_out0;
assign v_G22_1899_out0 = v_G11_13439_out0 && v_STALL_DUAL_CORE_4695_out0;
assign v_NOTUSED_1968_out0 = v__4856_out0;
assign v_NOTUSED_1969_out0 = v__4857_out0;
assign v_SIG_RD_11bit_3301_out0 = v__7714_out0;
assign v_SIG_RD_11bit_3302_out0 = v__7715_out0;
assign v_SIG_RM_11bit_6892_out0 = v__2771_out0;
assign v_SIG_RM_11bit_6893_out0 = v__2772_out0;
assign v_STALL_dual_core_8741_out0 = v_STALL_DUAL_CORE_1958_out0;
assign v_D1_8843_out0 = (v_AD3_10483_out0 == 2'b00) ? v_WEN3_1691_out0 : 1'h0;
assign v_D1_8843_out1 = (v_AD3_10483_out0 == 2'b01) ? v_WEN3_1691_out0 : 1'h0;
assign v_D1_8843_out2 = (v_AD3_10483_out0 == 2'b10) ? v_WEN3_1691_out0 : 1'h0;
assign v_D1_8843_out3 = (v_AD3_10483_out0 == 2'b11) ? v_WEN3_1691_out0 : 1'h0;
assign v__9805_out0 = { v__1952_out0,v_G3_207_out0 };
assign v__9807_out0 = { v__1954_out0,v_G3_209_out0 };
assign v__10262_out0 = { v_MUX13_13647_out0,v_0_10706_out0 };
assign v__10263_out0 = { v_MUX13_13648_out0,v_0_10707_out0 };
assign v__10370_out0 = { v_STALL_DUAL_CORE_4695_out0,v_C_1807_out0 };
assign v__10814_out0 = { v__4856_out1,v_C1_604_out0 };
assign v__10815_out0 = { v__4857_out1,v_C1_605_out0 };
assign v__10858_out0 = { v_MUX12_13783_out0,v_0_10706_out0 };
assign v__10859_out0 = { v_MUX12_13784_out0,v_0_10707_out0 };
assign v_OP2_SIG11_14_out0 = v_SIG_RM_11bit_6892_out0;
assign v_OP2_SIG11_15_out0 = v_SIG_RM_11bit_6893_out0;
assign v__73_out0 = { v__97_out0,v_G7_4822_out0 };
assign v_G4_219_out0 = v_G30_183_out0 || v_G3_2903_out0;
assign v_XOR3_2546_out0 = v_NEG1_6921_out0 ^ v__10858_out0;
assign v_XOR3_2547_out0 = v_NEG1_6922_out0 ^ v__10859_out0;
assign v_SUB_2909_out0 = v_G22_1899_out0;
assign v_MUX2_3255_out0 = v_LSR_6912_out0 ? v__10814_out0 : v_MUX1_31_out0;
assign v_MUX2_3256_out0 = v_LSR_6913_out0 ? v__10815_out0 : v_MUX1_32_out0;
assign v_EN_7093_out0 = v_STALL_dual_core_8741_out0;
assign v__8688_out0 = { v__9805_out0,v_G4_10998_out0 };
assign v__8690_out0 = { v__9807_out0,v_G4_11000_out0 };
assign v_RD_SIG11_8854_out0 = v_SIG_RD_11bit_3301_out0;
assign v_RD_SIG11_8855_out0 = v_SIG_RD_11bit_3302_out0;
assign v_A_10821_out0 = v__10370_out0;
assign v__60_out0 = v_A_10821_out0[10:10];
assign v__171_out0 = v_A_10821_out0[7:7];
assign v__179_out0 = v_A_10821_out0[3:3];
assign v__287_out0 = v_A_10821_out0[2:2];
assign v__1875_out0 = v_A_10821_out0[11:11];
assign v__2022_out0 = v_A_10821_out0[5:5];
assign v__2268_out0 = v_A_10821_out0[8:8];
assign v__3123_out0 = v_A_10821_out0[1:1];
assign v__3252_out0 = { v__8688_out0,v_G5_10569_out0 };
assign v__3254_out0 = { v__8690_out0,v_G5_10571_out0 };
assign v__3270_out0 = v_A_10821_out0[4:4];
assign v_MUX8_4587_out0 = v_MULTI_INSTRUCTION_13308_out0 ? v__10858_out0 : v_XOR3_2546_out0;
assign v_MUX8_4588_out0 = v_MULTI_INSTRUCTION_13309_out0 ? v__10859_out0 : v_XOR3_2547_out0;
assign v_OP2_SIG11_4827_out0 = v_OP2_SIG11_14_out0;
assign v_OP2_SIG11_4828_out0 = v_OP2_SIG11_15_out0;
assign v_RD_SIG11_7132_out0 = v_RD_SIG11_8854_out0;
assign v_RD_SIG11_7133_out0 = v_RD_SIG11_8855_out0;
assign v__8682_out0 = { v__73_out0,v_G8_2025_out0 };
assign v_Q_10339_out0 = v_OP2_SIG11_14_out0;
assign v_Q_10340_out0 = v_RD_SIG11_8854_out0;
assign v_Q_10341_out0 = v_OP2_SIG11_15_out0;
assign v_Q_10342_out0 = v_RD_SIG11_8855_out0;
assign v__11242_out0 = v_A_10821_out0[9:9];
assign v_IN_13306_out0 = v_MUX2_3255_out0;
assign v_IN_13307_out0 = v_MUX2_3256_out0;
assign v__13396_out0 = v_A_10821_out0[6:6];
assign v__13562_out0 = v_A_10821_out0[0:0];
assign v_WENLDST_13755_out0 = v_G4_219_out0;
assign v_G5_229_out0 = ((v__3270_out0 && !v_SUB_2909_out0) || (!v__3270_out0) && v_SUB_2909_out0);
assign v_G8_2024_out0 = ((v__171_out0 && !v_SUB_2909_out0) || (!v__171_out0) && v_SUB_2909_out0);
assign v_G9_2332_out0 = ((v__2268_out0 && !v_SUB_2909_out0) || (!v__2268_out0) && v_SUB_2909_out0);
assign v_G6_2416_out0 = ((v__2022_out0 && !v_SUB_2909_out0) || (!v__2022_out0) && v_SUB_2909_out0);
assign v_G11_2550_out0 = ((v__60_out0 && !v_SUB_2909_out0) || (!v__60_out0) && v_SUB_2909_out0);
assign v_G3_2621_out0 = ((v__287_out0 && !v_SUB_2909_out0) || (!v__287_out0) && v_SUB_2909_out0);
assign v_G10_2632_out0 = ((v__11242_out0 && !v_SUB_2909_out0) || (!v__11242_out0) && v_SUB_2909_out0);
assign v_WENLDST_2682_out0 = v_WENLDST_13755_out0;
assign v__2839_out0 = { v__8682_out0,v_G9_2333_out0 };
assign v__2889_out0 = v_IN_13306_out0[0:0];
assign v__2889_out1 = v_IN_13306_out0[15:15];
assign v__2890_out0 = v_IN_13307_out0[0:0];
assign v__2890_out1 = v_IN_13307_out0[15:15];
assign v_G2_3239_out0 = ((v__3123_out0 && !v_SUB_2909_out0) || (!v__3123_out0) && v_SUB_2909_out0);
assign v_G12_4699_out0 = ((v__1875_out0 && !v_SUB_2909_out0) || (!v__1875_out0) && v_SUB_2909_out0);
assign v_G7_4821_out0 = ((v__13396_out0 && !v_SUB_2909_out0) || (!v__13396_out0) && v_SUB_2909_out0);
assign v__7638_out0 = { v_Q_10339_out0,v_C1_10313_out0 };
assign v__7639_out0 = { v_Q_10340_out0,v_C1_10314_out0 };
assign v__7640_out0 = { v_Q_10341_out0,v_C1_10315_out0 };
assign v__7641_out0 = { v_Q_10342_out0,v_C1_10316_out0 };
assign v__10299_out0 = { v__3252_out0,v_G6_13638_out0 };
assign v__10301_out0 = { v__3254_out0,v_G6_13640_out0 };
assign v_G1_10477_out0 = ((v__13562_out0 && !v_SUB_2909_out0) || (!v__13562_out0) && v_SUB_2909_out0);
assign v__10808_out0 = v_IN_13306_out0[15:15];
assign v__10809_out0 = v_IN_13307_out0[15:15];
assign v_G4_12238_out0 = ((v__179_out0 && !v_SUB_2909_out0) || (!v__179_out0) && v_SUB_2909_out0);
assign {v_A4_13603_out1,v_A4_13603_out0 } = v__10262_out0 + v_MUX8_4587_out0 + v_G4_13702_out0;
assign {v_A4_13604_out1,v_A4_13604_out0 } = v__10263_out0 + v_MUX8_4588_out0 + v_G4_13703_out0;
assign v__120_out0 = { v__10299_out0,v_G7_2780_out0 };
assign v__122_out0 = { v__10301_out0,v_G7_2782_out0 };
assign v__333_out0 = { v__2889_out1,v__10808_out0 };
assign v__334_out0 = { v__2890_out1,v__10809_out0 };
assign v_WENLS_600_out0 = v_WENLDST_2682_out0;
assign v__1707_out0 = { v_G1_10477_out0,v_G2_3239_out0 };
assign v__2650_out0 = { v__2839_out0,v_G10_2633_out0 };
assign v_UNUSED1_3016_out0 = v_A4_13603_out1;
assign v_UNUSED1_3017_out0 = v_A4_13604_out1;
assign v_NOTUSED_4463_out0 = v__2889_out0;
assign v_NOTUSED_4464_out0 = v__2890_out0;
assign v_EXP_SUM_5844_out0 = v_A4_13603_out0;
assign v_EXP_SUM_5845_out0 = v_A4_13604_out0;
assign v_OUT_7708_out0 = v__7638_out0;
assign v_OUT_7709_out0 = v__7639_out0;
assign v_OUT_7710_out0 = v__7640_out0;
assign v_OUT_7711_out0 = v__7641_out0;
assign v_MUX3_8817_out0 = v_IR15_2464_out0 ? v_WENALU_8659_out0 : v_WENLDST_2682_out0;
assign v_SEL2_10323_out0 = v_A4_13603_out0[5:5];
assign v_SEL2_10324_out0 = v_A4_13604_out0[5:5];
assign v_RD_MULTI_45_out0 = v_OUT_7709_out0;
assign v_RD_MULTI_46_out0 = v_OUT_7711_out0;
assign v_RM_MULTI_210_out0 = v_OUT_7708_out0;
assign v_RM_MULTI_211_out0 = v_OUT_7710_out0;
assign v__2386_out0 = { v__1707_out0,v_G3_2621_out0 };
assign {v_A6_3957_out1,v_A6_3957_out0 } = v_EXP_SUM_5844_out0 + v_MUX10_10395_out0 + v_0_10706_out0;
assign {v_A6_3958_out1,v_A6_3958_out0 } = v_EXP_SUM_5845_out0 + v_MUX10_10396_out0 + v_0_10707_out0;
assign v__4734_out0 = { v__2650_out0,v_G11_2551_out0 };
assign v_XOR4_6960_out0 = v_EXP_SUM_5844_out0 ^ v_NEG1_6921_out0;
assign v_XOR4_6961_out0 = v_EXP_SUM_5845_out0 ^ v_NEG1_6922_out0;
assign v_MUX6_8757_out0 = v_MULTI_OPCODE_3020_out0 ? v_WEN_MULTI_2388_out0 : v_MUX3_8817_out0;
assign v_OUT_11234_out0 = v__333_out0;
assign v_OUT_11235_out0 = v__334_out0;
assign v_NEGATIVE_11256_out0 = v_SEL2_10323_out0;
assign v_NEGATIVE_11257_out0 = v_SEL2_10324_out0;
assign v_WENLS_11260_out0 = v_WENLS_600_out0;
assign v__13791_out0 = { v__120_out0,v_G8_1216_out0 };
assign v__13793_out0 = { v__122_out0,v_G8_1218_out0 };
assign v_WWNELS1_47_out0 = v_WENLS_11260_out0;
assign v_MUX4_275_out0 = v_NEGATIVE_11256_out0 ? v_OP2_EXP_10383_out0 : v_RD_EXP_2601_out0;
assign v_MUX4_276_out0 = v_NEGATIVE_11257_out0 ? v_OP2_EXP_10384_out0 : v_RD_EXP_2602_out0;
assign v__465_out0 = { v__13791_out0,v_G9_13286_out0 };
assign v__467_out0 = { v__13793_out0,v_G9_13288_out0 };
assign v_RM_MULTI_648_out0 = v_RM_MULTI_210_out0;
assign v_RM_MULTI_649_out0 = v_RM_MULTI_211_out0;
assign v_WEN3_1690_out0 = v_MUX6_8757_out0;
assign v_UNUSED2_2193_out0 = v_A6_3957_out1;
assign v_UNUSED2_2194_out0 = v_A6_3958_out1;
assign v_SHIFT_RD_2544_out0 = v_NEGATIVE_11256_out0;
assign v_SHIFT_RD_2545_out0 = v_NEGATIVE_11257_out0;
assign {v_A5_2638_out1,v_A5_2638_out0 } = v_XOR4_6960_out0 + v_C11_13765_out0 + v_C10_1819_out0;
assign {v_A5_2639_out1,v_A5_2639_out0 } = v_XOR4_6961_out0 + v_C11_13766_out0 + v_C10_1820_out0;
assign v_RD_FLOATING_2823_out0 = v_RD_MULTI_45_out0;
assign v_RD_FLOATING_2824_out0 = v_RD_MULTI_46_out0;
assign v__2968_out0 = { v__2386_out0,v_G4_12238_out0 };
assign v_SEL4_5790_out0 = v_A6_3957_out0[4:0];
assign v_SEL4_5791_out0 = v_A6_3958_out0[4:0];
assign v_MUX3_7075_out0 = v_ASR_8754_out0 ? v_OUT_11234_out0 : v_MUX2_3255_out0;
assign v_MUX3_7076_out0 = v_ASR_8755_out0 ? v_OUT_11235_out0 : v_MUX2_3256_out0;
assign v__10784_out0 = { v__4734_out0,v_G12_4700_out0 };
assign v_MUX11_86_out0 = v_G5_7106_out0 ? v_SEL4_5790_out0 : v_MUX4_275_out0;
assign v_MUX11_87_out0 = v_G5_7107_out0 ? v_SEL4_5791_out0 : v_MUX4_276_out0;
assign v_UNUSED_339_out0 = v_A5_2638_out1;
assign v_UNUSED_340_out0 = v_A5_2639_out1;
assign v__423_out0 = { v__465_out0,v_G10_13216_out0 };
assign v__425_out0 = { v__467_out0,v_G10_13218_out0 };
assign v_MUX7_1165_out0 = v_FLOATING_INS_13797_out0 ? v_RD_FLOATING_2823_out0 : v_RD_501_out0;
assign v_MUX7_1166_out0 = v_FLOATING_INS_13798_out0 ? v_RD_FLOATING_2824_out0 : v_RD_502_out0;
assign v_MUX8_1907_out0 = v_FLOATING_INS_13797_out0 ? v_RM_MULTI_648_out0 : v_RM_13750_out0;
assign v_MUX8_1908_out0 = v_FLOATING_INS_13798_out0 ? v_RM_MULTI_649_out0 : v_RM_13751_out0;
assign v__2984_out0 = v_MUX3_7075_out0[0:0];
assign v__2984_out1 = v_MUX3_7075_out0[15:15];
assign v__2985_out0 = v_MUX3_7076_out0[0:0];
assign v__2985_out1 = v_MUX3_7076_out0[15:15];
assign v__5849_out0 = { v__2968_out0,v_G5_229_out0 };
assign v_D1_8842_out0 = (v_AD3_10482_out0 == 2'b00) ? v_WEN3_1690_out0 : 1'h0;
assign v_D1_8842_out1 = (v_AD3_10482_out0 == 2'b01) ? v_WEN3_1690_out0 : 1'h0;
assign v_D1_8842_out2 = (v_AD3_10482_out0 == 2'b10) ? v_WEN3_1690_out0 : 1'h0;
assign v_D1_8842_out3 = (v_AD3_10482_out0 == 2'b11) ? v_WEN3_1690_out0 : 1'h0;
assign v_G1_10757_out0 = ! v_SHIFT_RD_2544_out0;
assign v_G1_10758_out0 = ! v_SHIFT_RD_2545_out0;
assign v_ADDER_IN_10996_out0 = v__10784_out0;
assign v_MUX9_13486_out0 = v_NEGATIVE_11256_out0 ? v_A5_2638_out0 : v_EXP_SUM_5844_out0;
assign v_MUX9_13487_out0 = v_NEGATIVE_11257_out0 ? v_A5_2639_out0 : v_EXP_SUM_5845_out0;
assign v__96_out0 = { v__5849_out0,v_G6_2416_out0 };
assign v_SEL3_390_out0 = v_MUX9_13486_out0[4:0];
assign v_SEL3_391_out0 = v_MUX9_13487_out0[4:0];
assign v_RD_613_out0 = v_MUX7_1165_out0;
assign v_RD_614_out0 = v_MUX7_1166_out0;
assign v__2835_out0 = { v__423_out0,v_G11_13343_out0 };
assign v__2837_out0 = { v__425_out0,v_G11_13345_out0 };
assign v_RM_3272_out0 = v_MUX8_1907_out0;
assign v_RM_3273_out0 = v_MUX8_1908_out0;
assign v__7120_out0 = { v__2984_out1,v__2984_out0 };
assign v__7121_out0 = { v__2985_out1,v__2985_out0 };
assign v_SHIFT_WHICH_OP_10715_out0 = v_G1_10757_out0;
assign v_SHIFT_WHICH_OP_10716_out0 = v_G1_10758_out0;
assign v_EXP_ANS_10860_out0 = v_MUX11_86_out0;
assign v_EXP_ANS_10861_out0 = v_MUX11_87_out0;
assign v__72_out0 = { v__96_out0,v_G7_4821_out0 };
assign v__437_out0 = v_RD_613_out0[2:2];
assign v__438_out0 = v_RD_614_out0[2:2];
assign v__2692_out0 = v_RD_613_out0[1:1];
assign v__2693_out0 = v_RD_614_out0[1:1];
assign v_RM_2912_out0 = v_RM_3272_out0;
assign v_RM_2913_out0 = v_RM_3273_out0;
assign v__3180_out0 = v_RD_613_out0[3:3];
assign v__3181_out0 = v_RD_614_out0[3:3];
assign v_SHIFT_WHICH_OP_4459_out0 = v_SHIFT_WHICH_OP_10715_out0;
assign v_SHIFT_WHICH_OP_4460_out0 = v_SHIFT_WHICH_OP_10716_out0;
assign v_SHIFT_AMOUNT_4715_out0 = v_SEL3_390_out0;
assign v_SHIFT_AMOUNT_4716_out0 = v_SEL3_391_out0;
assign v_RD_4839_out0 = v_RD_613_out0;
assign v_RD_4840_out0 = v_RD_614_out0;
assign v_MUX4_7023_out0 = v_ROR_3288_out0 ? v__7120_out0 : v_MUX3_7075_out0;
assign v_MUX4_7024_out0 = v_ROR_3289_out0 ? v__7121_out0 : v_MUX3_7076_out0;
assign v__7108_out0 = v_RD_613_out0[0:0];
assign v__7109_out0 = v_RD_614_out0[0:0];
assign v_A_10274_out0 = v_RM_3272_out0;
assign v_A_10276_out0 = v_RM_3273_out0;
assign v_SHIFT_WHICH_OP_10465_out0 = v_SHIFT_WHICH_OP_10715_out0;
assign v_SHIFT_WHICH_OP_10466_out0 = v_SHIFT_WHICH_OP_10716_out0;
assign v_EXP_PRE_ANS_10765_out0 = v_EXP_ANS_10860_out0;
assign v_EXP_PRE_ANS_10766_out0 = v_EXP_ANS_10861_out0;
assign v_RM_11064_out0 = v_RM_3272_out0;
assign v_RM_11065_out0 = v_RM_3272_out0;
assign v_RM_11067_out0 = v_RM_3272_out0;
assign v_RM_11079_out0 = v_RM_3273_out0;
assign v_RM_11080_out0 = v_RM_3273_out0;
assign v_RM_11082_out0 = v_RM_3273_out0;
assign v__11138_out0 = { v__2835_out0,v_G12_3346_out0 };
assign v__11140_out0 = { v__2837_out0,v_G12_3348_out0 };
assign v__0_out0 = v_A_10274_out0[4:4];
assign v__2_out0 = v_A_10276_out0[4:4];
assign v__37_out0 = v_RD_4839_out0[7:7];
assign v__38_out0 = v_RD_4840_out0[7:7];
assign v_SHIFT_AMOUNT_226_out0 = v_SHIFT_AMOUNT_4715_out0;
assign v_SHIFT_AMOUNT_227_out0 = v_SHIFT_AMOUNT_4716_out0;
assign v__504_out0 = v_RM_11064_out0[5:5];
assign v__505_out0 = v_RM_11065_out0[5:5];
assign v__507_out0 = v_RM_11067_out0[5:5];
assign v__519_out0 = v_RM_11079_out0[5:5];
assign v__520_out0 = v_RM_11080_out0[5:5];
assign v__522_out0 = v_RM_11082_out0[5:5];
assign v__569_out0 = v_RM_11064_out0[1:1];
assign v__570_out0 = v_RM_11065_out0[1:1];
assign v__572_out0 = v_RM_11067_out0[1:1];
assign v__584_out0 = v_RM_11079_out0[1:1];
assign v__585_out0 = v_RM_11080_out0[1:1];
assign v__587_out0 = v_RM_11082_out0[1:1];
assign v__1176_out0 = v_RD_4839_out0[13:13];
assign v__1177_out0 = v_RD_4840_out0[13:13];
assign v__1193_out0 = v_RD_4839_out0[4:4];
assign v__1194_out0 = v_RD_4840_out0[4:4];
assign v__1692_out0 = v_A_10274_out0[5:5];
assign v__1694_out0 = v_A_10276_out0[5:5];
assign v__1747_out0 = v_A_10274_out0[11:11];
assign v__1749_out0 = v_A_10276_out0[11:11];
assign v__1893_out0 = v_A_10274_out0[0:0];
assign v__1895_out0 = v_A_10276_out0[0:0];
assign v__1976_out0 = v_RM_11064_out0[15:15];
assign v__1977_out0 = v_RM_11065_out0[15:15];
assign v__1979_out0 = v_RM_11067_out0[15:15];
assign v__1991_out0 = v_RM_11079_out0[15:15];
assign v__1992_out0 = v_RM_11080_out0[15:15];
assign v__1994_out0 = v_RM_11082_out0[15:15];
assign v__2064_out0 = v_RM_11064_out0[10:10];
assign v__2065_out0 = v_RM_11065_out0[10:10];
assign v__2067_out0 = v_RM_11067_out0[10:10];
assign v__2079_out0 = v_RM_11079_out0[10:10];
assign v__2080_out0 = v_RM_11080_out0[10:10];
assign v__2082_out0 = v_RM_11082_out0[10:10];
assign v__2150_out0 = v_A_10274_out0[2:2];
assign v__2152_out0 = v_A_10276_out0[2:2];
assign v__2274_out0 = v_RM_11064_out0[12:12];
assign v__2275_out0 = v_RM_11065_out0[12:12];
assign v__2277_out0 = v_RM_11067_out0[12:12];
assign v__2289_out0 = v_RM_11079_out0[12:12];
assign v__2290_out0 = v_RM_11080_out0[12:12];
assign v__2292_out0 = v_RM_11082_out0[12:12];
assign v_MUX1_2401_out0 = v_SHIFT_WHICH_OP_10465_out0 ? v__2771_out0 : v__7714_out0;
assign v_MUX1_2402_out0 = v_SHIFT_WHICH_OP_10466_out0 ? v__2772_out0 : v__7715_out0;
assign v__2467_out0 = v_RD_4839_out0[8:8];
assign v__2468_out0 = v_RD_4840_out0[8:8];
assign v__2727_out0 = v_RM_11064_out0[2:2];
assign v__2728_out0 = v_RM_11065_out0[2:2];
assign v__2730_out0 = v_RM_11067_out0[2:2];
assign v__2742_out0 = v_RM_11079_out0[2:2];
assign v__2743_out0 = v_RM_11080_out0[2:2];
assign v__2745_out0 = v_RM_11082_out0[2:2];
assign v__2760_out0 = v_A_10274_out0[15:15];
assign v__2762_out0 = v_A_10276_out0[15:15];
assign v__2875_out0 = v_A_10274_out0[12:12];
assign v__2877_out0 = v_A_10276_out0[12:12];
assign v__2879_out0 = v_A_10274_out0[3:3];
assign v__2881_out0 = v_A_10276_out0[3:3];
assign v_EXP_2907_out0 = v_EXP_PRE_ANS_10765_out0;
assign v_EXP_2908_out0 = v_EXP_PRE_ANS_10766_out0;
assign v__2973_out0 = v_RD_4839_out0[15:15];
assign v__2974_out0 = v_RD_4840_out0[15:15];
assign v__2987_out0 = v_RM_11064_out0[8:8];
assign v__2988_out0 = v_RM_11065_out0[8:8];
assign v__2990_out0 = v_RM_11067_out0[8:8];
assign v__3002_out0 = v_RM_11079_out0[8:8];
assign v__3003_out0 = v_RM_11080_out0[8:8];
assign v__3005_out0 = v_RM_11082_out0[8:8];
assign v__3193_out0 = { v__11138_out0,v_G13_4706_out0 };
assign v__3195_out0 = { v__11140_out0,v_G13_4708_out0 };
assign v__3199_out0 = v_RD_4839_out0[10:10];
assign v__3200_out0 = v_RD_4840_out0[10:10];
assign v__3247_out0 = v_A_10274_out0[8:8];
assign v__3249_out0 = v_A_10276_out0[8:8];
assign v_RDN_3349_out0 = v__7108_out0;
assign v_RDN_3351_out0 = v__7109_out0;
assign v__3803_out0 = v_RD_4839_out0[12:12];
assign v__3804_out0 = v_RD_4840_out0[12:12];
assign v__3911_out0 = v_RM_11064_out0[11:11];
assign v__3912_out0 = v_RM_11065_out0[11:11];
assign v__3914_out0 = v_RM_11067_out0[11:11];
assign v__3926_out0 = v_RM_11079_out0[11:11];
assign v__3927_out0 = v_RM_11080_out0[11:11];
assign v__3929_out0 = v_RM_11082_out0[11:11];
assign v__3962_out0 = v_RM_11064_out0[9:9];
assign v__3963_out0 = v_RM_11065_out0[9:9];
assign v__3965_out0 = v_RM_11067_out0[9:9];
assign v__3977_out0 = v_RM_11079_out0[9:9];
assign v__3978_out0 = v_RM_11080_out0[9:9];
assign v__3980_out0 = v_RM_11082_out0[9:9];
assign v_RDN_4497_out0 = v__2692_out0;
assign v_RDN_4498_out0 = v__437_out0;
assign v_RDN_4500_out0 = v__3180_out0;
assign v_RDN_4512_out0 = v__2693_out0;
assign v_RDN_4513_out0 = v__438_out0;
assign v_RDN_4515_out0 = v__3181_out0;
assign v__4597_out0 = v_A_10274_out0[10:10];
assign v__4599_out0 = v_A_10276_out0[10:10];
assign v__4711_out0 = v_A_10274_out0[13:13];
assign v__4713_out0 = v_A_10276_out0[13:13];
assign v__6831_out0 = v_RM_11064_out0[14:14];
assign v__6832_out0 = v_RM_11065_out0[14:14];
assign v__6834_out0 = v_RM_11067_out0[14:14];
assign v__6846_out0 = v_RM_11079_out0[14:14];
assign v__6847_out0 = v_RM_11080_out0[14:14];
assign v__6849_out0 = v_RM_11082_out0[14:14];
assign v_MUX5_7017_out0 = v_EN_2330_out0 ? v_MUX4_7023_out0 : v_IN_13788_out0;
assign v_MUX5_7018_out0 = v_EN_2331_out0 ? v_MUX4_7024_out0 : v_IN_13789_out0;
assign v__8681_out0 = { v__72_out0,v_G8_2024_out0 };
assign v__8848_out0 = v_A_10274_out0[14:14];
assign v__8850_out0 = v_A_10276_out0[14:14];
assign v__10410_out0 = v_RM_11064_out0[7:7];
assign v__10411_out0 = v_RM_11065_out0[7:7];
assign v__10413_out0 = v_RM_11067_out0[7:7];
assign v__10425_out0 = v_RM_11079_out0[7:7];
assign v__10426_out0 = v_RM_11080_out0[7:7];
assign v__10428_out0 = v_RM_11082_out0[7:7];
assign v__10472_out0 = v_RD_4839_out0[9:9];
assign v__10473_out0 = v_RD_4840_out0[9:9];
assign v__10479_out0 = v_RD_4839_out0[6:6];
assign v__10480_out0 = v_RD_4840_out0[6:6];
assign v__10717_out0 = v_RD_4839_out0[14:14];
assign v__10718_out0 = v_RD_4840_out0[14:14];
assign v__10875_out0 = v_RM_11064_out0[4:4];
assign v__10876_out0 = v_RM_11065_out0[4:4];
assign v__10878_out0 = v_RM_11067_out0[4:4];
assign v__10890_out0 = v_RM_11079_out0[4:4];
assign v__10891_out0 = v_RM_11080_out0[4:4];
assign v__10893_out0 = v_RM_11082_out0[4:4];
assign v__11002_out0 = v_RM_11064_out0[0:0];
assign v__11003_out0 = v_RM_11065_out0[0:0];
assign v__11005_out0 = v_RM_11067_out0[0:0];
assign v__11017_out0 = v_RM_11079_out0[0:0];
assign v__11018_out0 = v_RM_11080_out0[0:0];
assign v__11020_out0 = v_RM_11082_out0[0:0];
assign v_RM_11063_out0 = v_RM_2912_out0;
assign v_RM_11066_out0 = v_RM_2912_out0;
assign v_RM_11068_out0 = v_RM_2912_out0;
assign v_RM_11069_out0 = v_RM_2912_out0;
assign v_RM_11070_out0 = v_RM_2912_out0;
assign v_RM_11071_out0 = v_RM_2912_out0;
assign v_RM_11072_out0 = v_RM_2912_out0;
assign v_RM_11073_out0 = v_RM_2912_out0;
assign v_RM_11074_out0 = v_RM_2912_out0;
assign v_RM_11075_out0 = v_RM_2912_out0;
assign v_RM_11076_out0 = v_RM_2912_out0;
assign v_RM_11077_out0 = v_RM_2912_out0;
assign v_RM_11078_out0 = v_RM_2913_out0;
assign v_RM_11081_out0 = v_RM_2913_out0;
assign v_RM_11083_out0 = v_RM_2913_out0;
assign v_RM_11084_out0 = v_RM_2913_out0;
assign v_RM_11085_out0 = v_RM_2913_out0;
assign v_RM_11086_out0 = v_RM_2913_out0;
assign v_RM_11087_out0 = v_RM_2913_out0;
assign v_RM_11088_out0 = v_RM_2913_out0;
assign v_RM_11089_out0 = v_RM_2913_out0;
assign v_RM_11090_out0 = v_RM_2913_out0;
assign v_RM_11091_out0 = v_RM_2913_out0;
assign v_RM_11092_out0 = v_RM_2913_out0;
assign v__11099_out0 = v_RM_11064_out0[3:3];
assign v__11100_out0 = v_RM_11065_out0[3:3];
assign v__11102_out0 = v_RM_11067_out0[3:3];
assign v__11114_out0 = v_RM_11079_out0[3:3];
assign v__11115_out0 = v_RM_11080_out0[3:3];
assign v__11117_out0 = v_RM_11082_out0[3:3];
assign v__11149_out0 = v_A_10274_out0[6:6];
assign v__11151_out0 = v_A_10276_out0[6:6];
assign v__13384_out0 = v_A_10274_out0[7:7];
assign v__13386_out0 = v_A_10276_out0[7:7];
assign v__13400_out0 = v_RM_11064_out0[6:6];
assign v__13401_out0 = v_RM_11065_out0[6:6];
assign v__13403_out0 = v_RM_11067_out0[6:6];
assign v__13415_out0 = v_RM_11079_out0[6:6];
assign v__13416_out0 = v_RM_11080_out0[6:6];
assign v__13418_out0 = v_RM_11082_out0[6:6];
assign v__13435_out0 = v_RD_4839_out0[5:5];
assign v__13436_out0 = v_RD_4840_out0[5:5];
assign v__13512_out0 = v_A_10274_out0[1:1];
assign v__13514_out0 = v_A_10276_out0[1:1];
assign v__13601_out0 = v_RD_4839_out0[11:11];
assign v__13602_out0 = v_RD_4840_out0[11:11];
assign v__13627_out0 = v_A_10274_out0[9:9];
assign v__13629_out0 = v_A_10276_out0[9:9];
assign v__13716_out0 = v_RM_11064_out0[13:13];
assign v__13717_out0 = v_RM_11065_out0[13:13];
assign v__13719_out0 = v_RM_11067_out0[13:13];
assign v__13731_out0 = v_RM_11079_out0[13:13];
assign v__13732_out0 = v_RM_11080_out0[13:13];
assign v__13734_out0 = v_RM_11082_out0[13:13];
assign v__174_out0 = { v__3193_out0,v_G14_4534_out0 };
assign v__176_out0 = { v__3195_out0,v_G14_4536_out0 };
assign v_G3_242_out0 = v_RDN_4497_out0 && v__2727_out0;
assign v_G3_243_out0 = v_RDN_4498_out0 && v__2728_out0;
assign v_G3_245_out0 = v_RDN_4500_out0 && v__2730_out0;
assign v_G3_257_out0 = v_RDN_4512_out0 && v__2742_out0;
assign v_G3_258_out0 = v_RDN_4513_out0 && v__2743_out0;
assign v_G3_260_out0 = v_RDN_4515_out0 && v__2745_out0;
assign v_G4_342_out0 = v_RDN_4497_out0 && v__11099_out0;
assign v_G4_343_out0 = v_RDN_4498_out0 && v__11100_out0;
assign v_G4_345_out0 = v_RDN_4500_out0 && v__11102_out0;
assign v_G4_357_out0 = v_RDN_4512_out0 && v__11114_out0;
assign v_G4_358_out0 = v_RDN_4513_out0 && v__11115_out0;
assign v_G4_360_out0 = v_RDN_4515_out0 && v__11117_out0;
assign v__503_out0 = v_RM_11063_out0[5:5];
assign v__506_out0 = v_RM_11066_out0[5:5];
assign v__508_out0 = v_RM_11068_out0[5:5];
assign v__509_out0 = v_RM_11069_out0[5:5];
assign v__510_out0 = v_RM_11070_out0[5:5];
assign v__511_out0 = v_RM_11071_out0[5:5];
assign v__512_out0 = v_RM_11072_out0[5:5];
assign v__513_out0 = v_RM_11073_out0[5:5];
assign v__514_out0 = v_RM_11074_out0[5:5];
assign v__515_out0 = v_RM_11075_out0[5:5];
assign v__516_out0 = v_RM_11076_out0[5:5];
assign v__517_out0 = v_RM_11077_out0[5:5];
assign v__518_out0 = v_RM_11078_out0[5:5];
assign v__521_out0 = v_RM_11081_out0[5:5];
assign v__523_out0 = v_RM_11083_out0[5:5];
assign v__524_out0 = v_RM_11084_out0[5:5];
assign v__525_out0 = v_RM_11085_out0[5:5];
assign v__526_out0 = v_RM_11086_out0[5:5];
assign v__527_out0 = v_RM_11087_out0[5:5];
assign v__528_out0 = v_RM_11088_out0[5:5];
assign v__529_out0 = v_RM_11089_out0[5:5];
assign v__530_out0 = v_RM_11090_out0[5:5];
assign v__531_out0 = v_RM_11091_out0[5:5];
assign v__532_out0 = v_RM_11092_out0[5:5];
assign v_G8_548_out0 = v__13384_out0 && v_RDN_3349_out0;
assign v_G8_550_out0 = v__13386_out0 && v_RDN_3351_out0;
assign v__568_out0 = v_RM_11063_out0[1:1];
assign v__571_out0 = v_RM_11066_out0[1:1];
assign v__573_out0 = v_RM_11068_out0[1:1];
assign v__574_out0 = v_RM_11069_out0[1:1];
assign v__575_out0 = v_RM_11070_out0[1:1];
assign v__576_out0 = v_RM_11071_out0[1:1];
assign v__577_out0 = v_RM_11072_out0[1:1];
assign v__578_out0 = v_RM_11073_out0[1:1];
assign v__579_out0 = v_RM_11074_out0[1:1];
assign v__580_out0 = v_RM_11075_out0[1:1];
assign v__581_out0 = v_RM_11076_out0[1:1];
assign v__582_out0 = v_RM_11077_out0[1:1];
assign v__583_out0 = v_RM_11078_out0[1:1];
assign v__586_out0 = v_RM_11081_out0[1:1];
assign v__588_out0 = v_RM_11083_out0[1:1];
assign v__589_out0 = v_RM_11084_out0[1:1];
assign v__590_out0 = v_RM_11085_out0[1:1];
assign v__591_out0 = v_RM_11086_out0[1:1];
assign v__592_out0 = v_RM_11087_out0[1:1];
assign v__593_out0 = v_RM_11088_out0[1:1];
assign v__594_out0 = v_RM_11089_out0[1:1];
assign v__595_out0 = v_RM_11090_out0[1:1];
assign v__596_out0 = v_RM_11091_out0[1:1];
assign v__597_out0 = v_RM_11092_out0[1:1];
assign v_G14_615_out0 = v__4711_out0 && v_RDN_3349_out0;
assign v_G14_617_out0 = v__4713_out0 && v_RDN_3351_out0;
assign v_G13_642_out0 = v__2875_out0 && v_RDN_3349_out0;
assign v_G13_644_out0 = v__2877_out0 && v_RDN_3351_out0;
assign v_OUT_1136_out0 = v_MUX5_7017_out0;
assign v_OUT_1137_out0 = v_MUX5_7018_out0;
assign v_G2_1809_out0 = v__13512_out0 && v_RDN_3349_out0;
assign v_G2_1811_out0 = v__13514_out0 && v_RDN_3351_out0;
assign v_G1_1879_out0 = v__1893_out0 && v_RDN_3349_out0;
assign v_G1_1881_out0 = v__1895_out0 && v_RDN_3351_out0;
assign v_G1_1910_out0 = v_RDN_4497_out0 && v__569_out0;
assign v_G1_1911_out0 = v_RDN_4498_out0 && v__570_out0;
assign v_G1_1913_out0 = v_RDN_4500_out0 && v__572_out0;
assign v_G1_1925_out0 = v_RDN_4512_out0 && v__584_out0;
assign v_G1_1926_out0 = v_RDN_4513_out0 && v__585_out0;
assign v_G1_1928_out0 = v_RDN_4515_out0 && v__587_out0;
assign v__1975_out0 = v_RM_11063_out0[15:15];
assign v__1978_out0 = v_RM_11066_out0[15:15];
assign v__1980_out0 = v_RM_11068_out0[15:15];
assign v__1981_out0 = v_RM_11069_out0[15:15];
assign v__1982_out0 = v_RM_11070_out0[15:15];
assign v__1983_out0 = v_RM_11071_out0[15:15];
assign v__1984_out0 = v_RM_11072_out0[15:15];
assign v__1985_out0 = v_RM_11073_out0[15:15];
assign v__1986_out0 = v_RM_11074_out0[15:15];
assign v__1987_out0 = v_RM_11075_out0[15:15];
assign v__1988_out0 = v_RM_11076_out0[15:15];
assign v__1989_out0 = v_RM_11077_out0[15:15];
assign v__1990_out0 = v_RM_11078_out0[15:15];
assign v__1993_out0 = v_RM_11081_out0[15:15];
assign v__1995_out0 = v_RM_11083_out0[15:15];
assign v__1996_out0 = v_RM_11084_out0[15:15];
assign v__1997_out0 = v_RM_11085_out0[15:15];
assign v__1998_out0 = v_RM_11086_out0[15:15];
assign v__1999_out0 = v_RM_11087_out0[15:15];
assign v__2000_out0 = v_RM_11088_out0[15:15];
assign v__2001_out0 = v_RM_11089_out0[15:15];
assign v__2002_out0 = v_RM_11090_out0[15:15];
assign v__2003_out0 = v_RM_11091_out0[15:15];
assign v__2004_out0 = v_RM_11092_out0[15:15];
assign v__2063_out0 = v_RM_11063_out0[10:10];
assign v__2066_out0 = v_RM_11066_out0[10:10];
assign v__2068_out0 = v_RM_11068_out0[10:10];
assign v__2069_out0 = v_RM_11069_out0[10:10];
assign v__2070_out0 = v_RM_11070_out0[10:10];
assign v__2071_out0 = v_RM_11071_out0[10:10];
assign v__2072_out0 = v_RM_11072_out0[10:10];
assign v__2073_out0 = v_RM_11073_out0[10:10];
assign v__2074_out0 = v_RM_11074_out0[10:10];
assign v__2075_out0 = v_RM_11075_out0[10:10];
assign v__2076_out0 = v_RM_11076_out0[10:10];
assign v__2077_out0 = v_RM_11077_out0[10:10];
assign v__2078_out0 = v_RM_11078_out0[10:10];
assign v__2081_out0 = v_RM_11081_out0[10:10];
assign v__2083_out0 = v_RM_11083_out0[10:10];
assign v__2084_out0 = v_RM_11084_out0[10:10];
assign v__2085_out0 = v_RM_11085_out0[10:10];
assign v__2086_out0 = v_RM_11086_out0[10:10];
assign v__2087_out0 = v_RM_11087_out0[10:10];
assign v__2088_out0 = v_RM_11088_out0[10:10];
assign v__2089_out0 = v_RM_11089_out0[10:10];
assign v__2090_out0 = v_RM_11090_out0[10:10];
assign v__2091_out0 = v_RM_11091_out0[10:10];
assign v__2092_out0 = v_RM_11092_out0[10:10];
assign v_G6_2117_out0 = v_RDN_4497_out0 && v__13400_out0;
assign v_G6_2118_out0 = v_RDN_4498_out0 && v__13401_out0;
assign v_G6_2120_out0 = v_RDN_4500_out0 && v__13403_out0;
assign v_G6_2132_out0 = v_RDN_4512_out0 && v__13415_out0;
assign v_G6_2133_out0 = v_RDN_4513_out0 && v__13416_out0;
assign v_G6_2135_out0 = v_RDN_4515_out0 && v__13418_out0;
assign v__2273_out0 = v_RM_11063_out0[12:12];
assign v__2276_out0 = v_RM_11066_out0[12:12];
assign v__2278_out0 = v_RM_11068_out0[12:12];
assign v__2279_out0 = v_RM_11069_out0[12:12];
assign v__2280_out0 = v_RM_11070_out0[12:12];
assign v__2281_out0 = v_RM_11071_out0[12:12];
assign v__2282_out0 = v_RM_11072_out0[12:12];
assign v__2283_out0 = v_RM_11073_out0[12:12];
assign v__2284_out0 = v_RM_11074_out0[12:12];
assign v__2285_out0 = v_RM_11075_out0[12:12];
assign v__2286_out0 = v_RM_11076_out0[12:12];
assign v__2287_out0 = v_RM_11077_out0[12:12];
assign v__2288_out0 = v_RM_11078_out0[12:12];
assign v__2291_out0 = v_RM_11081_out0[12:12];
assign v__2293_out0 = v_RM_11083_out0[12:12];
assign v__2294_out0 = v_RM_11084_out0[12:12];
assign v__2295_out0 = v_RM_11085_out0[12:12];
assign v__2296_out0 = v_RM_11086_out0[12:12];
assign v__2297_out0 = v_RM_11087_out0[12:12];
assign v__2298_out0 = v_RM_11088_out0[12:12];
assign v__2299_out0 = v_RM_11089_out0[12:12];
assign v__2300_out0 = v_RM_11090_out0[12:12];
assign v__2301_out0 = v_RM_11091_out0[12:12];
assign v__2302_out0 = v_RM_11092_out0[12:12];
assign v_EXP_2441_out0 = v_EXP_2907_out0;
assign v_EXP_2442_out0 = v_EXP_2908_out0;
assign v_G8_2473_out0 = v_RDN_4497_out0 && v__2987_out0;
assign v_G8_2474_out0 = v_RDN_4498_out0 && v__2988_out0;
assign v_G8_2476_out0 = v_RDN_4500_out0 && v__2990_out0;
assign v_G8_2488_out0 = v_RDN_4512_out0 && v__3002_out0;
assign v_G8_2489_out0 = v_RDN_4513_out0 && v__3003_out0;
assign v_G8_2491_out0 = v_RDN_4515_out0 && v__3005_out0;
assign v_G10_2640_out0 = v__13627_out0 && v_RDN_3349_out0;
assign v_G10_2642_out0 = v__13629_out0 && v_RDN_3351_out0;
assign v__2726_out0 = v_RM_11063_out0[2:2];
assign v__2729_out0 = v_RM_11066_out0[2:2];
assign v__2731_out0 = v_RM_11068_out0[2:2];
assign v__2732_out0 = v_RM_11069_out0[2:2];
assign v__2733_out0 = v_RM_11070_out0[2:2];
assign v__2734_out0 = v_RM_11071_out0[2:2];
assign v__2735_out0 = v_RM_11072_out0[2:2];
assign v__2736_out0 = v_RM_11073_out0[2:2];
assign v__2737_out0 = v_RM_11074_out0[2:2];
assign v__2738_out0 = v_RM_11075_out0[2:2];
assign v__2739_out0 = v_RM_11076_out0[2:2];
assign v__2740_out0 = v_RM_11077_out0[2:2];
assign v__2741_out0 = v_RM_11078_out0[2:2];
assign v__2744_out0 = v_RM_11081_out0[2:2];
assign v__2746_out0 = v_RM_11083_out0[2:2];
assign v__2747_out0 = v_RM_11084_out0[2:2];
assign v__2748_out0 = v_RM_11085_out0[2:2];
assign v__2749_out0 = v_RM_11086_out0[2:2];
assign v__2750_out0 = v_RM_11087_out0[2:2];
assign v__2751_out0 = v_RM_11088_out0[2:2];
assign v__2752_out0 = v_RM_11089_out0[2:2];
assign v__2753_out0 = v_RM_11090_out0[2:2];
assign v__2754_out0 = v_RM_11091_out0[2:2];
assign v__2755_out0 = v_RM_11092_out0[2:2];
assign v_G4_2767_out0 = v__2879_out0 && v_RDN_3349_out0;
assign v_G4_2769_out0 = v__2881_out0 && v_RDN_3351_out0;
assign v_G5_2783_out0 = v__0_out0 && v_RDN_3349_out0;
assign v_G5_2785_out0 = v__2_out0 && v_RDN_3351_out0;
assign v__2838_out0 = { v__8681_out0,v_G9_2332_out0 };
assign v_G9_2895_out0 = v__3247_out0 && v_RDN_3349_out0;
assign v_G9_2897_out0 = v__3249_out0 && v_RDN_3351_out0;
assign v_G11_2937_out0 = v__4597_out0 && v_RDN_3349_out0;
assign v_G11_2939_out0 = v__4599_out0 && v_RDN_3351_out0;
assign v__2986_out0 = v_RM_11063_out0[8:8];
assign v__2989_out0 = v_RM_11066_out0[8:8];
assign v__2991_out0 = v_RM_11068_out0[8:8];
assign v__2992_out0 = v_RM_11069_out0[8:8];
assign v__2993_out0 = v_RM_11070_out0[8:8];
assign v__2994_out0 = v_RM_11071_out0[8:8];
assign v__2995_out0 = v_RM_11072_out0[8:8];
assign v__2996_out0 = v_RM_11073_out0[8:8];
assign v__2997_out0 = v_RM_11074_out0[8:8];
assign v__2998_out0 = v_RM_11075_out0[8:8];
assign v__2999_out0 = v_RM_11076_out0[8:8];
assign v__3000_out0 = v_RM_11077_out0[8:8];
assign v__3001_out0 = v_RM_11078_out0[8:8];
assign v__3004_out0 = v_RM_11081_out0[8:8];
assign v__3006_out0 = v_RM_11083_out0[8:8];
assign v__3007_out0 = v_RM_11084_out0[8:8];
assign v__3008_out0 = v_RM_11085_out0[8:8];
assign v__3009_out0 = v_RM_11086_out0[8:8];
assign v__3010_out0 = v_RM_11087_out0[8:8];
assign v__3011_out0 = v_RM_11088_out0[8:8];
assign v__3012_out0 = v_RM_11089_out0[8:8];
assign v__3013_out0 = v_RM_11090_out0[8:8];
assign v__3014_out0 = v_RM_11091_out0[8:8];
assign v__3015_out0 = v_RM_11092_out0[8:8];
assign v__3910_out0 = v_RM_11063_out0[11:11];
assign v__3913_out0 = v_RM_11066_out0[11:11];
assign v__3915_out0 = v_RM_11068_out0[11:11];
assign v__3916_out0 = v_RM_11069_out0[11:11];
assign v__3917_out0 = v_RM_11070_out0[11:11];
assign v__3918_out0 = v_RM_11071_out0[11:11];
assign v__3919_out0 = v_RM_11072_out0[11:11];
assign v__3920_out0 = v_RM_11073_out0[11:11];
assign v__3921_out0 = v_RM_11074_out0[11:11];
assign v__3922_out0 = v_RM_11075_out0[11:11];
assign v__3923_out0 = v_RM_11076_out0[11:11];
assign v__3924_out0 = v_RM_11077_out0[11:11];
assign v__3925_out0 = v_RM_11078_out0[11:11];
assign v__3928_out0 = v_RM_11081_out0[11:11];
assign v__3930_out0 = v_RM_11083_out0[11:11];
assign v__3931_out0 = v_RM_11084_out0[11:11];
assign v__3932_out0 = v_RM_11085_out0[11:11];
assign v__3933_out0 = v_RM_11086_out0[11:11];
assign v__3934_out0 = v_RM_11087_out0[11:11];
assign v__3935_out0 = v_RM_11088_out0[11:11];
assign v__3936_out0 = v_RM_11089_out0[11:11];
assign v__3937_out0 = v_RM_11090_out0[11:11];
assign v__3938_out0 = v_RM_11091_out0[11:11];
assign v__3939_out0 = v_RM_11092_out0[11:11];
assign v_B_3946_out0 = v_SHIFT_AMOUNT_226_out0;
assign v_B_3947_out0 = v_SHIFT_AMOUNT_227_out0;
assign v__3961_out0 = v_RM_11063_out0[9:9];
assign v__3964_out0 = v_RM_11066_out0[9:9];
assign v__3966_out0 = v_RM_11068_out0[9:9];
assign v__3967_out0 = v_RM_11069_out0[9:9];
assign v__3968_out0 = v_RM_11070_out0[9:9];
assign v__3969_out0 = v_RM_11071_out0[9:9];
assign v__3970_out0 = v_RM_11072_out0[9:9];
assign v__3971_out0 = v_RM_11073_out0[9:9];
assign v__3972_out0 = v_RM_11074_out0[9:9];
assign v__3973_out0 = v_RM_11075_out0[9:9];
assign v__3974_out0 = v_RM_11076_out0[9:9];
assign v__3975_out0 = v_RM_11077_out0[9:9];
assign v__3976_out0 = v_RM_11078_out0[9:9];
assign v__3979_out0 = v_RM_11081_out0[9:9];
assign v__3981_out0 = v_RM_11083_out0[9:9];
assign v__3982_out0 = v_RM_11084_out0[9:9];
assign v__3983_out0 = v_RM_11085_out0[9:9];
assign v__3984_out0 = v_RM_11086_out0[9:9];
assign v__3985_out0 = v_RM_11087_out0[9:9];
assign v__3986_out0 = v_RM_11088_out0[9:9];
assign v__3987_out0 = v_RM_11089_out0[9:9];
assign v__3988_out0 = v_RM_11090_out0[9:9];
assign v__3989_out0 = v_RM_11091_out0[9:9];
assign v__3990_out0 = v_RM_11092_out0[9:9];
assign v_RDN_4496_out0 = v__1193_out0;
assign v_RDN_4499_out0 = v__13601_out0;
assign v_RDN_4501_out0 = v__3199_out0;
assign v_RDN_4502_out0 = v__2973_out0;
assign v_RDN_4503_out0 = v__10717_out0;
assign v_RDN_4504_out0 = v__3803_out0;
assign v_RDN_4505_out0 = v__2467_out0;
assign v_RDN_4506_out0 = v__13435_out0;
assign v_RDN_4507_out0 = v__37_out0;
assign v_RDN_4508_out0 = v__1176_out0;
assign v_RDN_4509_out0 = v__10479_out0;
assign v_RDN_4510_out0 = v__10472_out0;
assign v_RDN_4511_out0 = v__1194_out0;
assign v_RDN_4514_out0 = v__13602_out0;
assign v_RDN_4516_out0 = v__3200_out0;
assign v_RDN_4517_out0 = v__2974_out0;
assign v_RDN_4518_out0 = v__10718_out0;
assign v_RDN_4519_out0 = v__3804_out0;
assign v_RDN_4520_out0 = v__2468_out0;
assign v_RDN_4521_out0 = v__13436_out0;
assign v_RDN_4522_out0 = v__38_out0;
assign v_RDN_4523_out0 = v__1177_out0;
assign v_RDN_4524_out0 = v__10480_out0;
assign v_RDN_4525_out0 = v__10473_out0;
assign v_G2_4621_out0 = v_RDN_4497_out0 && v__10875_out0;
assign v_G2_4622_out0 = v_RDN_4498_out0 && v__10876_out0;
assign v_G2_4624_out0 = v_RDN_4500_out0 && v__10878_out0;
assign v_G2_4636_out0 = v_RDN_4512_out0 && v__10890_out0;
assign v_G2_4637_out0 = v_RDN_4513_out0 && v__10891_out0;
assign v_G2_4639_out0 = v_RDN_4515_out0 && v__10893_out0;
assign v_G15_4654_out0 = v__8848_out0 && v_RDN_3349_out0;
assign v_G15_4656_out0 = v__8850_out0 && v_RDN_3351_out0;
assign v__6830_out0 = v_RM_11063_out0[14:14];
assign v__6833_out0 = v_RM_11066_out0[14:14];
assign v__6835_out0 = v_RM_11068_out0[14:14];
assign v__6836_out0 = v_RM_11069_out0[14:14];
assign v__6837_out0 = v_RM_11070_out0[14:14];
assign v__6838_out0 = v_RM_11071_out0[14:14];
assign v__6839_out0 = v_RM_11072_out0[14:14];
assign v__6840_out0 = v_RM_11073_out0[14:14];
assign v__6841_out0 = v_RM_11074_out0[14:14];
assign v__6842_out0 = v_RM_11075_out0[14:14];
assign v__6843_out0 = v_RM_11076_out0[14:14];
assign v__6844_out0 = v_RM_11077_out0[14:14];
assign v__6845_out0 = v_RM_11078_out0[14:14];
assign v__6848_out0 = v_RM_11081_out0[14:14];
assign v__6850_out0 = v_RM_11083_out0[14:14];
assign v__6851_out0 = v_RM_11084_out0[14:14];
assign v__6852_out0 = v_RM_11085_out0[14:14];
assign v__6853_out0 = v_RM_11086_out0[14:14];
assign v__6854_out0 = v_RM_11087_out0[14:14];
assign v__6855_out0 = v_RM_11088_out0[14:14];
assign v__6856_out0 = v_RM_11089_out0[14:14];
assign v__6857_out0 = v_RM_11090_out0[14:14];
assign v__6858_out0 = v_RM_11091_out0[14:14];
assign v__6859_out0 = v_RM_11092_out0[14:14];
assign v_EQ1_6956_out0 = v_EXP_2907_out0 == 5'h0;
assign v_EQ1_6957_out0 = v_EXP_2908_out0 == 5'h0;
assign v_G3_7087_out0 = v__2150_out0 && v_RDN_3349_out0;
assign v_G3_7089_out0 = v__2152_out0 && v_RDN_3351_out0;
assign v_G7_8655_out0 = v__11149_out0 && v_RDN_3349_out0;
assign v_G7_8657_out0 = v__11151_out0 && v_RDN_3351_out0;
assign v_G6_8834_out0 = v__1692_out0 && v_RDN_3349_out0;
assign v_G6_8836_out0 = v__1694_out0 && v_RDN_3351_out0;
assign v__10409_out0 = v_RM_11063_out0[7:7];
assign v__10412_out0 = v_RM_11066_out0[7:7];
assign v__10414_out0 = v_RM_11068_out0[7:7];
assign v__10415_out0 = v_RM_11069_out0[7:7];
assign v__10416_out0 = v_RM_11070_out0[7:7];
assign v__10417_out0 = v_RM_11071_out0[7:7];
assign v__10418_out0 = v_RM_11072_out0[7:7];
assign v__10419_out0 = v_RM_11073_out0[7:7];
assign v__10420_out0 = v_RM_11074_out0[7:7];
assign v__10421_out0 = v_RM_11075_out0[7:7];
assign v__10422_out0 = v_RM_11076_out0[7:7];
assign v__10423_out0 = v_RM_11077_out0[7:7];
assign v__10424_out0 = v_RM_11078_out0[7:7];
assign v__10427_out0 = v_RM_11081_out0[7:7];
assign v__10429_out0 = v_RM_11083_out0[7:7];
assign v__10430_out0 = v_RM_11084_out0[7:7];
assign v__10431_out0 = v_RM_11085_out0[7:7];
assign v__10432_out0 = v_RM_11086_out0[7:7];
assign v__10433_out0 = v_RM_11087_out0[7:7];
assign v__10434_out0 = v_RM_11088_out0[7:7];
assign v__10435_out0 = v_RM_11089_out0[7:7];
assign v__10436_out0 = v_RM_11090_out0[7:7];
assign v__10437_out0 = v_RM_11091_out0[7:7];
assign v__10438_out0 = v_RM_11092_out0[7:7];
assign v_G9_10573_out0 = v_RDN_4497_out0 && v__3962_out0;
assign v_G9_10574_out0 = v_RDN_4498_out0 && v__3963_out0;
assign v_G9_10576_out0 = v_RDN_4500_out0 && v__3965_out0;
assign v_G9_10588_out0 = v_RDN_4512_out0 && v__3977_out0;
assign v_G9_10589_out0 = v_RDN_4513_out0 && v__3978_out0;
assign v_G9_10591_out0 = v_RDN_4515_out0 && v__3980_out0;
assign v_G5_10622_out0 = v_RDN_4497_out0 && v__504_out0;
assign v_G5_10623_out0 = v_RDN_4498_out0 && v__505_out0;
assign v_G5_10625_out0 = v_RDN_4500_out0 && v__507_out0;
assign v_G5_10637_out0 = v_RDN_4512_out0 && v__519_out0;
assign v_G5_10638_out0 = v_RDN_4513_out0 && v__520_out0;
assign v_G5_10640_out0 = v_RDN_4515_out0 && v__522_out0;
assign v_G12_10688_out0 = v__1747_out0 && v_RDN_3349_out0;
assign v_G12_10690_out0 = v__1749_out0 && v_RDN_3351_out0;
assign v_SIG_TO_SHIFT_10712_out0 = v_MUX1_2401_out0;
assign v_SIG_TO_SHIFT_10713_out0 = v_MUX1_2402_out0;
assign v__10874_out0 = v_RM_11063_out0[4:4];
assign v__10877_out0 = v_RM_11066_out0[4:4];
assign v__10879_out0 = v_RM_11068_out0[4:4];
assign v__10880_out0 = v_RM_11069_out0[4:4];
assign v__10881_out0 = v_RM_11070_out0[4:4];
assign v__10882_out0 = v_RM_11071_out0[4:4];
assign v__10883_out0 = v_RM_11072_out0[4:4];
assign v__10884_out0 = v_RM_11073_out0[4:4];
assign v__10885_out0 = v_RM_11074_out0[4:4];
assign v__10886_out0 = v_RM_11075_out0[4:4];
assign v__10887_out0 = v_RM_11076_out0[4:4];
assign v__10888_out0 = v_RM_11077_out0[4:4];
assign v__10889_out0 = v_RM_11078_out0[4:4];
assign v__10892_out0 = v_RM_11081_out0[4:4];
assign v__10894_out0 = v_RM_11083_out0[4:4];
assign v__10895_out0 = v_RM_11084_out0[4:4];
assign v__10896_out0 = v_RM_11085_out0[4:4];
assign v__10897_out0 = v_RM_11086_out0[4:4];
assign v__10898_out0 = v_RM_11087_out0[4:4];
assign v__10899_out0 = v_RM_11088_out0[4:4];
assign v__10900_out0 = v_RM_11089_out0[4:4];
assign v__10901_out0 = v_RM_11090_out0[4:4];
assign v__10902_out0 = v_RM_11091_out0[4:4];
assign v__10903_out0 = v_RM_11092_out0[4:4];
assign v_G16_10906_out0 = v__2760_out0 && v_RDN_3349_out0;
assign v_G16_10908_out0 = v__2762_out0 && v_RDN_3351_out0;
assign v__11001_out0 = v_RM_11063_out0[0:0];
assign v__11004_out0 = v_RM_11066_out0[0:0];
assign v__11006_out0 = v_RM_11068_out0[0:0];
assign v__11007_out0 = v_RM_11069_out0[0:0];
assign v__11008_out0 = v_RM_11070_out0[0:0];
assign v__11009_out0 = v_RM_11071_out0[0:0];
assign v__11010_out0 = v_RM_11072_out0[0:0];
assign v__11011_out0 = v_RM_11073_out0[0:0];
assign v__11012_out0 = v_RM_11074_out0[0:0];
assign v__11013_out0 = v_RM_11075_out0[0:0];
assign v__11014_out0 = v_RM_11076_out0[0:0];
assign v__11015_out0 = v_RM_11077_out0[0:0];
assign v__11016_out0 = v_RM_11078_out0[0:0];
assign v__11019_out0 = v_RM_11081_out0[0:0];
assign v__11021_out0 = v_RM_11083_out0[0:0];
assign v__11022_out0 = v_RM_11084_out0[0:0];
assign v__11023_out0 = v_RM_11085_out0[0:0];
assign v__11024_out0 = v_RM_11086_out0[0:0];
assign v__11025_out0 = v_RM_11087_out0[0:0];
assign v__11026_out0 = v_RM_11088_out0[0:0];
assign v__11027_out0 = v_RM_11089_out0[0:0];
assign v__11028_out0 = v_RM_11090_out0[0:0];
assign v__11029_out0 = v_RM_11091_out0[0:0];
assign v__11030_out0 = v_RM_11092_out0[0:0];
assign v__11098_out0 = v_RM_11063_out0[3:3];
assign v__11101_out0 = v_RM_11066_out0[3:3];
assign v__11103_out0 = v_RM_11068_out0[3:3];
assign v__11104_out0 = v_RM_11069_out0[3:3];
assign v__11105_out0 = v_RM_11070_out0[3:3];
assign v__11106_out0 = v_RM_11071_out0[3:3];
assign v__11107_out0 = v_RM_11072_out0[3:3];
assign v__11108_out0 = v_RM_11073_out0[3:3];
assign v__11109_out0 = v_RM_11074_out0[3:3];
assign v__11110_out0 = v_RM_11075_out0[3:3];
assign v__11111_out0 = v_RM_11076_out0[3:3];
assign v__11112_out0 = v_RM_11077_out0[3:3];
assign v__11113_out0 = v_RM_11078_out0[3:3];
assign v__11116_out0 = v_RM_11081_out0[3:3];
assign v__11118_out0 = v_RM_11083_out0[3:3];
assign v__11119_out0 = v_RM_11084_out0[3:3];
assign v__11120_out0 = v_RM_11085_out0[3:3];
assign v__11121_out0 = v_RM_11086_out0[3:3];
assign v__11122_out0 = v_RM_11087_out0[3:3];
assign v__11123_out0 = v_RM_11088_out0[3:3];
assign v__11124_out0 = v_RM_11089_out0[3:3];
assign v__11125_out0 = v_RM_11090_out0[3:3];
assign v__11126_out0 = v_RM_11091_out0[3:3];
assign v__11127_out0 = v_RM_11092_out0[3:3];
assign v_EQ2_11254_out0 = v_EXP_2907_out0 == 5'h1;
assign v_EQ2_11255_out0 = v_EXP_2908_out0 == 5'h1;
assign v_G7_11263_out0 = v_RDN_4497_out0 && v__10410_out0;
assign v_G7_11264_out0 = v_RDN_4498_out0 && v__10411_out0;
assign v_G7_11266_out0 = v_RDN_4500_out0 && v__10413_out0;
assign v_G7_11278_out0 = v_RDN_4512_out0 && v__10425_out0;
assign v_G7_11279_out0 = v_RDN_4513_out0 && v__10426_out0;
assign v_G7_11281_out0 = v_RDN_4515_out0 && v__10428_out0;
assign v_G16_13184_out0 = v_RDN_4497_out0 && v__11002_out0;
assign v_G16_13185_out0 = v_RDN_4498_out0 && v__11003_out0;
assign v_G16_13187_out0 = v_RDN_4500_out0 && v__11005_out0;
assign v_G16_13199_out0 = v_RDN_4512_out0 && v__11017_out0;
assign v_G16_13200_out0 = v_RDN_4513_out0 && v__11018_out0;
assign v_G16_13202_out0 = v_RDN_4515_out0 && v__11020_out0;
assign v__13399_out0 = v_RM_11063_out0[6:6];
assign v__13402_out0 = v_RM_11066_out0[6:6];
assign v__13404_out0 = v_RM_11068_out0[6:6];
assign v__13405_out0 = v_RM_11069_out0[6:6];
assign v__13406_out0 = v_RM_11070_out0[6:6];
assign v__13407_out0 = v_RM_11071_out0[6:6];
assign v__13408_out0 = v_RM_11072_out0[6:6];
assign v__13409_out0 = v_RM_11073_out0[6:6];
assign v__13410_out0 = v_RM_11074_out0[6:6];
assign v__13411_out0 = v_RM_11075_out0[6:6];
assign v__13412_out0 = v_RM_11076_out0[6:6];
assign v__13413_out0 = v_RM_11077_out0[6:6];
assign v__13414_out0 = v_RM_11078_out0[6:6];
assign v__13417_out0 = v_RM_11081_out0[6:6];
assign v__13419_out0 = v_RM_11083_out0[6:6];
assign v__13420_out0 = v_RM_11084_out0[6:6];
assign v__13421_out0 = v_RM_11085_out0[6:6];
assign v__13422_out0 = v_RM_11086_out0[6:6];
assign v__13423_out0 = v_RM_11087_out0[6:6];
assign v__13424_out0 = v_RM_11088_out0[6:6];
assign v__13425_out0 = v_RM_11089_out0[6:6];
assign v__13426_out0 = v_RM_11090_out0[6:6];
assign v__13427_out0 = v_RM_11091_out0[6:6];
assign v__13428_out0 = v_RM_11092_out0[6:6];
assign v_RD_13568_out0 = v_RDN_4497_out0;
assign v_RD_13569_out0 = v_RDN_4498_out0;
assign v_RD_13571_out0 = v_RDN_4500_out0;
assign v_RD_13583_out0 = v_RDN_4512_out0;
assign v_RD_13584_out0 = v_RDN_4513_out0;
assign v_RD_13586_out0 = v_RDN_4515_out0;
assign v__13715_out0 = v_RM_11063_out0[13:13];
assign v__13718_out0 = v_RM_11066_out0[13:13];
assign v__13720_out0 = v_RM_11068_out0[13:13];
assign v__13721_out0 = v_RM_11069_out0[13:13];
assign v__13722_out0 = v_RM_11070_out0[13:13];
assign v__13723_out0 = v_RM_11071_out0[13:13];
assign v__13724_out0 = v_RM_11072_out0[13:13];
assign v__13725_out0 = v_RM_11073_out0[13:13];
assign v__13726_out0 = v_RM_11074_out0[13:13];
assign v__13727_out0 = v_RM_11075_out0[13:13];
assign v__13728_out0 = v_RM_11076_out0[13:13];
assign v__13729_out0 = v_RM_11077_out0[13:13];
assign v__13730_out0 = v_RM_11078_out0[13:13];
assign v__13733_out0 = v_RM_11081_out0[13:13];
assign v__13735_out0 = v_RM_11083_out0[13:13];
assign v__13736_out0 = v_RM_11084_out0[13:13];
assign v__13737_out0 = v_RM_11085_out0[13:13];
assign v__13738_out0 = v_RM_11086_out0[13:13];
assign v__13739_out0 = v_RM_11087_out0[13:13];
assign v__13740_out0 = v_RM_11088_out0[13:13];
assign v__13741_out0 = v_RM_11089_out0[13:13];
assign v__13742_out0 = v_RM_11090_out0[13:13];
assign v__13743_out0 = v_RM_11091_out0[13:13];
assign v__13744_out0 = v_RM_11092_out0[13:13];
assign v_G15_133_out0 = v_RD_13568_out0 && v__1976_out0;
assign v_G15_134_out0 = v_RD_13569_out0 && v__1977_out0;
assign v_G15_136_out0 = v_RD_13571_out0 && v__1979_out0;
assign v_G15_148_out0 = v_RD_13583_out0 && v__1991_out0;
assign v_G15_149_out0 = v_RD_13584_out0 && v__1992_out0;
assign v_G15_151_out0 = v_RD_13586_out0 && v__1994_out0;
assign v_G3_241_out0 = v_RDN_4496_out0 && v__2726_out0;
assign v_G3_244_out0 = v_RDN_4499_out0 && v__2729_out0;
assign v_G3_246_out0 = v_RDN_4501_out0 && v__2731_out0;
assign v_G3_247_out0 = v_RDN_4502_out0 && v__2732_out0;
assign v_G3_248_out0 = v_RDN_4503_out0 && v__2733_out0;
assign v_G3_249_out0 = v_RDN_4504_out0 && v__2734_out0;
assign v_G3_250_out0 = v_RDN_4505_out0 && v__2735_out0;
assign v_G3_251_out0 = v_RDN_4506_out0 && v__2736_out0;
assign v_G3_252_out0 = v_RDN_4507_out0 && v__2737_out0;
assign v_G3_253_out0 = v_RDN_4508_out0 && v__2738_out0;
assign v_G3_254_out0 = v_RDN_4509_out0 && v__2739_out0;
assign v_G3_255_out0 = v_RDN_4510_out0 && v__2740_out0;
assign v_G3_256_out0 = v_RDN_4511_out0 && v__2741_out0;
assign v_G3_259_out0 = v_RDN_4514_out0 && v__2744_out0;
assign v_G3_261_out0 = v_RDN_4516_out0 && v__2746_out0;
assign v_G3_262_out0 = v_RDN_4517_out0 && v__2747_out0;
assign v_G3_263_out0 = v_RDN_4518_out0 && v__2748_out0;
assign v_G3_264_out0 = v_RDN_4519_out0 && v__2749_out0;
assign v_G3_265_out0 = v_RDN_4520_out0 && v__2750_out0;
assign v_G3_266_out0 = v_RDN_4521_out0 && v__2751_out0;
assign v_G3_267_out0 = v_RDN_4522_out0 && v__2752_out0;
assign v_G3_268_out0 = v_RDN_4523_out0 && v__2753_out0;
assign v_G3_269_out0 = v_RDN_4524_out0 && v__2754_out0;
assign v_G3_270_out0 = v_RDN_4525_out0 && v__2755_out0;
assign v_G4_341_out0 = v_RDN_4496_out0 && v__11098_out0;
assign v_G4_344_out0 = v_RDN_4499_out0 && v__11101_out0;
assign v_G4_346_out0 = v_RDN_4501_out0 && v__11103_out0;
assign v_G4_347_out0 = v_RDN_4502_out0 && v__11104_out0;
assign v_G4_348_out0 = v_RDN_4503_out0 && v__11105_out0;
assign v_G4_349_out0 = v_RDN_4504_out0 && v__11106_out0;
assign v_G4_350_out0 = v_RDN_4505_out0 && v__11107_out0;
assign v_G4_351_out0 = v_RDN_4506_out0 && v__11108_out0;
assign v_G4_352_out0 = v_RDN_4507_out0 && v__11109_out0;
assign v_G4_353_out0 = v_RDN_4508_out0 && v__11110_out0;
assign v_G4_354_out0 = v_RDN_4509_out0 && v__11111_out0;
assign v_G4_355_out0 = v_RDN_4510_out0 && v__11112_out0;
assign v_G4_356_out0 = v_RDN_4511_out0 && v__11113_out0;
assign v_G4_359_out0 = v_RDN_4514_out0 && v__11116_out0;
assign v_G4_361_out0 = v_RDN_4516_out0 && v__11118_out0;
assign v_G4_362_out0 = v_RDN_4517_out0 && v__11119_out0;
assign v_G4_363_out0 = v_RDN_4518_out0 && v__11120_out0;
assign v_G4_364_out0 = v_RDN_4519_out0 && v__11121_out0;
assign v_G4_365_out0 = v_RDN_4520_out0 && v__11122_out0;
assign v_G4_366_out0 = v_RDN_4521_out0 && v__11123_out0;
assign v_G4_367_out0 = v_RDN_4522_out0 && v__11124_out0;
assign v_G4_368_out0 = v_RDN_4523_out0 && v__11125_out0;
assign v_G4_369_out0 = v_RDN_4524_out0 && v__11126_out0;
assign v_G4_370_out0 = v_RDN_4525_out0 && v__11127_out0;
assign v__386_out0 = { v_G5_2783_out0,v_G6_8834_out0 };
assign v__388_out0 = { v_G5_2785_out0,v_G6_8836_out0 };
assign v__399_out0 = { v_G9_2895_out0,v_G10_2640_out0 };
assign v__401_out0 = { v_G9_2897_out0,v_G10_2642_out0 };
assign v_G11_652_out0 = v_RD_13568_out0 && v__3911_out0;
assign v_G11_653_out0 = v_RD_13569_out0 && v__3912_out0;
assign v_G11_655_out0 = v_RD_13571_out0 && v__3914_out0;
assign v_G11_667_out0 = v_RD_13583_out0 && v__3926_out0;
assign v_G11_668_out0 = v_RD_13584_out0 && v__3927_out0;
assign v_G11_670_out0 = v_RD_13586_out0 && v__3929_out0;
assign v_2_1763_out0 = v_B_3946_out0[2:2];
assign v_2_1764_out0 = v_B_3947_out0[2:2];
assign v_G1_1909_out0 = v_RDN_4496_out0 && v__568_out0;
assign v_G1_1912_out0 = v_RDN_4499_out0 && v__571_out0;
assign v_G1_1914_out0 = v_RDN_4501_out0 && v__573_out0;
assign v_G1_1915_out0 = v_RDN_4502_out0 && v__574_out0;
assign v_G1_1916_out0 = v_RDN_4503_out0 && v__575_out0;
assign v_G1_1917_out0 = v_RDN_4504_out0 && v__576_out0;
assign v_G1_1918_out0 = v_RDN_4505_out0 && v__577_out0;
assign v_G1_1919_out0 = v_RDN_4506_out0 && v__578_out0;
assign v_G1_1920_out0 = v_RDN_4507_out0 && v__579_out0;
assign v_G1_1921_out0 = v_RDN_4508_out0 && v__580_out0;
assign v_G1_1922_out0 = v_RDN_4509_out0 && v__581_out0;
assign v_G1_1923_out0 = v_RDN_4510_out0 && v__582_out0;
assign v_G1_1924_out0 = v_RDN_4511_out0 && v__583_out0;
assign v_G1_1927_out0 = v_RDN_4514_out0 && v__586_out0;
assign v_G1_1929_out0 = v_RDN_4516_out0 && v__588_out0;
assign v_G1_1930_out0 = v_RDN_4517_out0 && v__589_out0;
assign v_G1_1931_out0 = v_RDN_4518_out0 && v__590_out0;
assign v_G1_1932_out0 = v_RDN_4519_out0 && v__591_out0;
assign v_G1_1933_out0 = v_RDN_4520_out0 && v__592_out0;
assign v_G1_1934_out0 = v_RDN_4521_out0 && v__593_out0;
assign v_G1_1935_out0 = v_RDN_4522_out0 && v__594_out0;
assign v_G1_1936_out0 = v_RDN_4523_out0 && v__595_out0;
assign v_G1_1937_out0 = v_RDN_4524_out0 && v__596_out0;
assign v_G1_1938_out0 = v_RDN_4525_out0 && v__597_out0;
assign v_G6_2116_out0 = v_RDN_4496_out0 && v__13399_out0;
assign v_G6_2119_out0 = v_RDN_4499_out0 && v__13402_out0;
assign v_G6_2121_out0 = v_RDN_4501_out0 && v__13404_out0;
assign v_G6_2122_out0 = v_RDN_4502_out0 && v__13405_out0;
assign v_G6_2123_out0 = v_RDN_4503_out0 && v__13406_out0;
assign v_G6_2124_out0 = v_RDN_4504_out0 && v__13407_out0;
assign v_G6_2125_out0 = v_RDN_4505_out0 && v__13408_out0;
assign v_G6_2126_out0 = v_RDN_4506_out0 && v__13409_out0;
assign v_G6_2127_out0 = v_RDN_4507_out0 && v__13410_out0;
assign v_G6_2128_out0 = v_RDN_4508_out0 && v__13411_out0;
assign v_G6_2129_out0 = v_RDN_4509_out0 && v__13412_out0;
assign v_G6_2130_out0 = v_RDN_4510_out0 && v__13413_out0;
assign v_G6_2131_out0 = v_RDN_4511_out0 && v__13414_out0;
assign v_G6_2134_out0 = v_RDN_4514_out0 && v__13417_out0;
assign v_G6_2136_out0 = v_RDN_4516_out0 && v__13419_out0;
assign v_G6_2137_out0 = v_RDN_4517_out0 && v__13420_out0;
assign v_G6_2138_out0 = v_RDN_4518_out0 && v__13421_out0;
assign v_G6_2139_out0 = v_RDN_4519_out0 && v__13422_out0;
assign v_G6_2140_out0 = v_RDN_4520_out0 && v__13423_out0;
assign v_G6_2141_out0 = v_RDN_4521_out0 && v__13424_out0;
assign v_G6_2142_out0 = v_RDN_4522_out0 && v__13425_out0;
assign v_G6_2143_out0 = v_RDN_4523_out0 && v__13426_out0;
assign v_G6_2144_out0 = v_RDN_4524_out0 && v__13427_out0;
assign v_G6_2145_out0 = v_RDN_4525_out0 && v__13428_out0;
assign v_G8_2472_out0 = v_RDN_4496_out0 && v__2986_out0;
assign v_G8_2475_out0 = v_RDN_4499_out0 && v__2989_out0;
assign v_G8_2477_out0 = v_RDN_4501_out0 && v__2991_out0;
assign v_G8_2478_out0 = v_RDN_4502_out0 && v__2992_out0;
assign v_G8_2479_out0 = v_RDN_4503_out0 && v__2993_out0;
assign v_G8_2480_out0 = v_RDN_4504_out0 && v__2994_out0;
assign v_G8_2481_out0 = v_RDN_4505_out0 && v__2995_out0;
assign v_G8_2482_out0 = v_RDN_4506_out0 && v__2996_out0;
assign v_G8_2483_out0 = v_RDN_4507_out0 && v__2997_out0;
assign v_G8_2484_out0 = v_RDN_4508_out0 && v__2998_out0;
assign v_G8_2485_out0 = v_RDN_4509_out0 && v__2999_out0;
assign v_G8_2486_out0 = v_RDN_4510_out0 && v__3000_out0;
assign v_G8_2487_out0 = v_RDN_4511_out0 && v__3001_out0;
assign v_G8_2490_out0 = v_RDN_4514_out0 && v__3004_out0;
assign v_G8_2492_out0 = v_RDN_4516_out0 && v__3006_out0;
assign v_G8_2493_out0 = v_RDN_4517_out0 && v__3007_out0;
assign v_G8_2494_out0 = v_RDN_4518_out0 && v__3008_out0;
assign v_G8_2495_out0 = v_RDN_4519_out0 && v__3009_out0;
assign v_G8_2496_out0 = v_RDN_4520_out0 && v__3010_out0;
assign v_G8_2497_out0 = v_RDN_4521_out0 && v__3011_out0;
assign v_G8_2498_out0 = v_RDN_4522_out0 && v__3012_out0;
assign v_G8_2499_out0 = v_RDN_4523_out0 && v__3013_out0;
assign v_G8_2500_out0 = v_RDN_4524_out0 && v__3014_out0;
assign v_G8_2501_out0 = v_RDN_4525_out0 && v__3015_out0;
assign v__2649_out0 = { v__2838_out0,v_G10_2632_out0 };
assign v__2945_out0 = { v_G15_4654_out0,v_G16_10906_out0 };
assign v__2947_out0 = { v_G15_4656_out0,v_G16_10908_out0 };
assign v_0_3022_out0 = v_B_3946_out0[0:0];
assign v_0_3023_out0 = v_B_3947_out0[0:0];
assign v__3215_out0 = { v_G1_1879_out0,v_G2_1809_out0 };
assign v__3217_out0 = { v_G1_1881_out0,v_G2_1811_out0 };
assign v__3278_out0 = { v_G3_7087_out0,v_G4_2767_out0 };
assign v__3280_out0 = { v_G3_7089_out0,v_G4_2769_out0 };
assign v_1_3817_out0 = v_B_3946_out0[1:1];
assign v_1_3818_out0 = v_B_3947_out0[1:1];
assign v_G2_4620_out0 = v_RDN_4496_out0 && v__10874_out0;
assign v_G2_4623_out0 = v_RDN_4499_out0 && v__10877_out0;
assign v_G2_4625_out0 = v_RDN_4501_out0 && v__10879_out0;
assign v_G2_4626_out0 = v_RDN_4502_out0 && v__10880_out0;
assign v_G2_4627_out0 = v_RDN_4503_out0 && v__10881_out0;
assign v_G2_4628_out0 = v_RDN_4504_out0 && v__10882_out0;
assign v_G2_4629_out0 = v_RDN_4505_out0 && v__10883_out0;
assign v_G2_4630_out0 = v_RDN_4506_out0 && v__10884_out0;
assign v_G2_4631_out0 = v_RDN_4507_out0 && v__10885_out0;
assign v_G2_4632_out0 = v_RDN_4508_out0 && v__10886_out0;
assign v_G2_4633_out0 = v_RDN_4509_out0 && v__10887_out0;
assign v_G2_4634_out0 = v_RDN_4510_out0 && v__10888_out0;
assign v_G2_4635_out0 = v_RDN_4511_out0 && v__10889_out0;
assign v_G2_4638_out0 = v_RDN_4514_out0 && v__10892_out0;
assign v_G2_4640_out0 = v_RDN_4516_out0 && v__10894_out0;
assign v_G2_4641_out0 = v_RDN_4517_out0 && v__10895_out0;
assign v_G2_4642_out0 = v_RDN_4518_out0 && v__10896_out0;
assign v_G2_4643_out0 = v_RDN_4519_out0 && v__10897_out0;
assign v_G2_4644_out0 = v_RDN_4520_out0 && v__10898_out0;
assign v_G2_4645_out0 = v_RDN_4521_out0 && v__10899_out0;
assign v_G2_4646_out0 = v_RDN_4522_out0 && v__10900_out0;
assign v_G2_4647_out0 = v_RDN_4523_out0 && v__10901_out0;
assign v_G2_4648_out0 = v_RDN_4524_out0 && v__10902_out0;
assign v_G2_4649_out0 = v_RDN_4525_out0 && v__10903_out0;
assign v_SIG_TO_SHIFT_5836_out0 = v_SIG_TO_SHIFT_10712_out0;
assign v_SIG_TO_SHIFT_5837_out0 = v_SIG_TO_SHIFT_10713_out0;
assign v_RD_5903_out0 = v_G16_13184_out0;
assign v_RD_5935_out0 = v_G16_13185_out0;
assign v_RD_5997_out0 = v_G16_13187_out0;
assign v_RD_6367_out0 = v_G16_13199_out0;
assign v_RD_6399_out0 = v_G16_13200_out0;
assign v_RD_6461_out0 = v_G16_13202_out0;
assign v_G10_6976_out0 = v_RD_13568_out0 && v__2064_out0;
assign v_G10_6977_out0 = v_RD_13569_out0 && v__2065_out0;
assign v_G10_6979_out0 = v_RD_13571_out0 && v__2067_out0;
assign v_G10_6991_out0 = v_RD_13583_out0 && v__2079_out0;
assign v_G10_6992_out0 = v_RD_13584_out0 && v__2080_out0;
assign v_G10_6994_out0 = v_RD_13586_out0 && v__2082_out0;
assign v__7135_out0 = { v_G13_642_out0,v_G14_615_out0 };
assign v__7137_out0 = { v_G13_644_out0,v_G14_617_out0 };
assign v_RD_7204_out0 = v_G5_10622_out0;
assign v_RD_7205_out0 = v_G2_4621_out0;
assign v_RD_7207_out0 = v_G9_10573_out0;
assign v_RD_7209_out0 = v_G1_1910_out0;
assign v_RD_7210_out0 = v_G4_342_out0;
assign v_RD_7211_out0 = v_G6_2117_out0;
assign v_RD_7212_out0 = v_G7_11263_out0;
assign v_RD_7214_out0 = v_G8_2473_out0;
assign v_RD_7215_out0 = v_G3_242_out0;
assign v_RD_7219_out0 = v_G5_10623_out0;
assign v_RD_7220_out0 = v_G2_4622_out0;
assign v_RD_7222_out0 = v_G9_10574_out0;
assign v_RD_7224_out0 = v_G1_1911_out0;
assign v_RD_7225_out0 = v_G4_343_out0;
assign v_RD_7226_out0 = v_G6_2118_out0;
assign v_RD_7227_out0 = v_G7_11264_out0;
assign v_RD_7229_out0 = v_G8_2474_out0;
assign v_RD_7230_out0 = v_G3_243_out0;
assign v_RD_7249_out0 = v_G5_10625_out0;
assign v_RD_7250_out0 = v_G2_4624_out0;
assign v_RD_7252_out0 = v_G9_10576_out0;
assign v_RD_7254_out0 = v_G1_1913_out0;
assign v_RD_7255_out0 = v_G4_345_out0;
assign v_RD_7256_out0 = v_G6_2120_out0;
assign v_RD_7257_out0 = v_G7_11266_out0;
assign v_RD_7259_out0 = v_G8_2476_out0;
assign v_RD_7260_out0 = v_G3_245_out0;
assign v_RD_7428_out0 = v_G5_10637_out0;
assign v_RD_7429_out0 = v_G2_4636_out0;
assign v_RD_7431_out0 = v_G9_10588_out0;
assign v_RD_7433_out0 = v_G1_1925_out0;
assign v_RD_7434_out0 = v_G4_357_out0;
assign v_RD_7435_out0 = v_G6_2132_out0;
assign v_RD_7436_out0 = v_G7_11278_out0;
assign v_RD_7438_out0 = v_G8_2488_out0;
assign v_RD_7439_out0 = v_G3_257_out0;
assign v_RD_7443_out0 = v_G5_10638_out0;
assign v_RD_7444_out0 = v_G2_4637_out0;
assign v_RD_7446_out0 = v_G9_10589_out0;
assign v_RD_7448_out0 = v_G1_1926_out0;
assign v_RD_7449_out0 = v_G4_358_out0;
assign v_RD_7450_out0 = v_G6_2133_out0;
assign v_RD_7451_out0 = v_G7_11279_out0;
assign v_RD_7453_out0 = v_G8_2489_out0;
assign v_RD_7454_out0 = v_G3_258_out0;
assign v_RD_7473_out0 = v_G5_10640_out0;
assign v_RD_7474_out0 = v_G2_4639_out0;
assign v_RD_7476_out0 = v_G9_10591_out0;
assign v_RD_7478_out0 = v_G1_1928_out0;
assign v_RD_7479_out0 = v_G4_360_out0;
assign v_RD_7480_out0 = v_G6_2135_out0;
assign v_RD_7481_out0 = v_G7_11281_out0;
assign v_RD_7483_out0 = v_G8_2491_out0;
assign v_RD_7484_out0 = v_G3_260_out0;
assign v_SUBNORMAL_8808_out0 = v_EQ1_6956_out0;
assign v_SUBNORMAL_8809_out0 = v_EQ1_6957_out0;
assign v_IN_10403_out0 = v_OUT_1136_out0;
assign v_IN_10404_out0 = v_OUT_1137_out0;
assign v__10456_out0 = { v__174_out0,v_G15_1815_out0 };
assign v__10458_out0 = { v__176_out0,v_G15_1817_out0 };
assign v_G9_10572_out0 = v_RDN_4496_out0 && v__3961_out0;
assign v_G9_10575_out0 = v_RDN_4499_out0 && v__3964_out0;
assign v_G9_10577_out0 = v_RDN_4501_out0 && v__3966_out0;
assign v_G9_10578_out0 = v_RDN_4502_out0 && v__3967_out0;
assign v_G9_10579_out0 = v_RDN_4503_out0 && v__3968_out0;
assign v_G9_10580_out0 = v_RDN_4504_out0 && v__3969_out0;
assign v_G9_10581_out0 = v_RDN_4505_out0 && v__3970_out0;
assign v_G9_10582_out0 = v_RDN_4506_out0 && v__3971_out0;
assign v_G9_10583_out0 = v_RDN_4507_out0 && v__3972_out0;
assign v_G9_10584_out0 = v_RDN_4508_out0 && v__3973_out0;
assign v_G9_10585_out0 = v_RDN_4509_out0 && v__3974_out0;
assign v_G9_10586_out0 = v_RDN_4510_out0 && v__3975_out0;
assign v_G9_10587_out0 = v_RDN_4511_out0 && v__3976_out0;
assign v_G9_10590_out0 = v_RDN_4514_out0 && v__3979_out0;
assign v_G9_10592_out0 = v_RDN_4516_out0 && v__3981_out0;
assign v_G9_10593_out0 = v_RDN_4517_out0 && v__3982_out0;
assign v_G9_10594_out0 = v_RDN_4518_out0 && v__3983_out0;
assign v_G9_10595_out0 = v_RDN_4519_out0 && v__3984_out0;
assign v_G9_10596_out0 = v_RDN_4520_out0 && v__3985_out0;
assign v_G9_10597_out0 = v_RDN_4521_out0 && v__3986_out0;
assign v_G9_10598_out0 = v_RDN_4522_out0 && v__3987_out0;
assign v_G9_10599_out0 = v_RDN_4523_out0 && v__3988_out0;
assign v_G9_10600_out0 = v_RDN_4524_out0 && v__3989_out0;
assign v_G9_10601_out0 = v_RDN_4525_out0 && v__3990_out0;
assign v_G5_10621_out0 = v_RDN_4496_out0 && v__503_out0;
assign v_G5_10624_out0 = v_RDN_4499_out0 && v__506_out0;
assign v_G5_10626_out0 = v_RDN_4501_out0 && v__508_out0;
assign v_G5_10627_out0 = v_RDN_4502_out0 && v__509_out0;
assign v_G5_10628_out0 = v_RDN_4503_out0 && v__510_out0;
assign v_G5_10629_out0 = v_RDN_4504_out0 && v__511_out0;
assign v_G5_10630_out0 = v_RDN_4505_out0 && v__512_out0;
assign v_G5_10631_out0 = v_RDN_4506_out0 && v__513_out0;
assign v_G5_10632_out0 = v_RDN_4507_out0 && v__514_out0;
assign v_G5_10633_out0 = v_RDN_4508_out0 && v__515_out0;
assign v_G5_10634_out0 = v_RDN_4509_out0 && v__516_out0;
assign v_G5_10635_out0 = v_RDN_4510_out0 && v__517_out0;
assign v_G5_10636_out0 = v_RDN_4511_out0 && v__518_out0;
assign v_G5_10639_out0 = v_RDN_4514_out0 && v__521_out0;
assign v_G5_10641_out0 = v_RDN_4516_out0 && v__523_out0;
assign v_G5_10642_out0 = v_RDN_4517_out0 && v__524_out0;
assign v_G5_10643_out0 = v_RDN_4518_out0 && v__525_out0;
assign v_G5_10644_out0 = v_RDN_4519_out0 && v__526_out0;
assign v_G5_10645_out0 = v_RDN_4520_out0 && v__527_out0;
assign v_G5_10646_out0 = v_RDN_4521_out0 && v__528_out0;
assign v_G5_10647_out0 = v_RDN_4522_out0 && v__529_out0;
assign v_G5_10648_out0 = v_RDN_4523_out0 && v__530_out0;
assign v_G5_10649_out0 = v_RDN_4524_out0 && v__531_out0;
assign v_G5_10650_out0 = v_RDN_4525_out0 && v__532_out0;
assign v_G7_11262_out0 = v_RDN_4496_out0 && v__10409_out0;
assign v_G7_11265_out0 = v_RDN_4499_out0 && v__10412_out0;
assign v_G7_11267_out0 = v_RDN_4501_out0 && v__10414_out0;
assign v_G7_11268_out0 = v_RDN_4502_out0 && v__10415_out0;
assign v_G7_11269_out0 = v_RDN_4503_out0 && v__10416_out0;
assign v_G7_11270_out0 = v_RDN_4504_out0 && v__10417_out0;
assign v_G7_11271_out0 = v_RDN_4505_out0 && v__10418_out0;
assign v_G7_11272_out0 = v_RDN_4506_out0 && v__10419_out0;
assign v_G7_11273_out0 = v_RDN_4507_out0 && v__10420_out0;
assign v_G7_11274_out0 = v_RDN_4508_out0 && v__10421_out0;
assign v_G7_11275_out0 = v_RDN_4509_out0 && v__10422_out0;
assign v_G7_11276_out0 = v_RDN_4510_out0 && v__10423_out0;
assign v_G7_11277_out0 = v_RDN_4511_out0 && v__10424_out0;
assign v_G7_11280_out0 = v_RDN_4514_out0 && v__10427_out0;
assign v_G7_11282_out0 = v_RDN_4516_out0 && v__10429_out0;
assign v_G7_11283_out0 = v_RDN_4517_out0 && v__10430_out0;
assign v_G7_11284_out0 = v_RDN_4518_out0 && v__10431_out0;
assign v_G7_11285_out0 = v_RDN_4519_out0 && v__10432_out0;
assign v_G7_11286_out0 = v_RDN_4520_out0 && v__10433_out0;
assign v_G7_11287_out0 = v_RDN_4521_out0 && v__10434_out0;
assign v_G7_11288_out0 = v_RDN_4522_out0 && v__10435_out0;
assign v_G7_11289_out0 = v_RDN_4523_out0 && v__10436_out0;
assign v_G7_11290_out0 = v_RDN_4524_out0 && v__10437_out0;
assign v_G7_11291_out0 = v_RDN_4525_out0 && v__10438_out0;
assign v_G16_13183_out0 = v_RDN_4496_out0 && v__11001_out0;
assign v_G16_13186_out0 = v_RDN_4499_out0 && v__11004_out0;
assign v_G16_13188_out0 = v_RDN_4501_out0 && v__11006_out0;
assign v_G16_13189_out0 = v_RDN_4502_out0 && v__11007_out0;
assign v_G16_13190_out0 = v_RDN_4503_out0 && v__11008_out0;
assign v_G16_13191_out0 = v_RDN_4504_out0 && v__11009_out0;
assign v_G16_13192_out0 = v_RDN_4505_out0 && v__11010_out0;
assign v_G16_13193_out0 = v_RDN_4506_out0 && v__11011_out0;
assign v_G16_13194_out0 = v_RDN_4507_out0 && v__11012_out0;
assign v_G16_13195_out0 = v_RDN_4508_out0 && v__11013_out0;
assign v_G16_13196_out0 = v_RDN_4509_out0 && v__11014_out0;
assign v_G16_13197_out0 = v_RDN_4510_out0 && v__11015_out0;
assign v_G16_13198_out0 = v_RDN_4511_out0 && v__11016_out0;
assign v_G16_13201_out0 = v_RDN_4514_out0 && v__11019_out0;
assign v_G16_13203_out0 = v_RDN_4516_out0 && v__11021_out0;
assign v_G16_13204_out0 = v_RDN_4517_out0 && v__11022_out0;
assign v_G16_13205_out0 = v_RDN_4518_out0 && v__11023_out0;
assign v_G16_13206_out0 = v_RDN_4519_out0 && v__11024_out0;
assign v_G16_13207_out0 = v_RDN_4520_out0 && v__11025_out0;
assign v_G16_13208_out0 = v_RDN_4521_out0 && v__11026_out0;
assign v_G16_13209_out0 = v_RDN_4522_out0 && v__11027_out0;
assign v_G16_13210_out0 = v_RDN_4523_out0 && v__11028_out0;
assign v_G16_13211_out0 = v_RDN_4524_out0 && v__11029_out0;
assign v_G16_13212_out0 = v_RDN_4525_out0 && v__11030_out0;
assign v_G12_13222_out0 = v_RD_13568_out0 && v__2274_out0;
assign v_G12_13223_out0 = v_RD_13569_out0 && v__2275_out0;
assign v_G12_13225_out0 = v_RD_13571_out0 && v__2277_out0;
assign v_G12_13237_out0 = v_RD_13583_out0 && v__2289_out0;
assign v_G12_13238_out0 = v_RD_13584_out0 && v__2290_out0;
assign v_G12_13240_out0 = v_RD_13586_out0 && v__2292_out0;
assign v__13261_out0 = { v_G11_2937_out0,v_G12_10688_out0 };
assign v__13263_out0 = { v_G11_2939_out0,v_G12_10690_out0 };
assign v_G13_13353_out0 = v_RD_13568_out0 && v__13716_out0;
assign v_G13_13354_out0 = v_RD_13569_out0 && v__13717_out0;
assign v_G13_13356_out0 = v_RD_13571_out0 && v__13719_out0;
assign v_G13_13368_out0 = v_RD_13583_out0 && v__13731_out0;
assign v_G13_13369_out0 = v_RD_13584_out0 && v__13732_out0;
assign v_G13_13371_out0 = v_RD_13586_out0 && v__13734_out0;
assign v_EXP1_13488_out0 = v_EQ2_11254_out0;
assign v_EXP1_13489_out0 = v_EQ2_11255_out0;
assign v_RD_13567_out0 = v_RDN_4496_out0;
assign v_RD_13570_out0 = v_RDN_4499_out0;
assign v_RD_13572_out0 = v_RDN_4501_out0;
assign v_RD_13573_out0 = v_RDN_4502_out0;
assign v_RD_13574_out0 = v_RDN_4503_out0;
assign v_RD_13575_out0 = v_RDN_4504_out0;
assign v_RD_13576_out0 = v_RDN_4505_out0;
assign v_RD_13577_out0 = v_RDN_4506_out0;
assign v_RD_13578_out0 = v_RDN_4507_out0;
assign v_RD_13579_out0 = v_RDN_4508_out0;
assign v_RD_13580_out0 = v_RDN_4509_out0;
assign v_RD_13581_out0 = v_RDN_4510_out0;
assign v_RD_13582_out0 = v_RDN_4511_out0;
assign v_RD_13585_out0 = v_RDN_4514_out0;
assign v_RD_13587_out0 = v_RDN_4516_out0;
assign v_RD_13588_out0 = v_RDN_4517_out0;
assign v_RD_13589_out0 = v_RDN_4518_out0;
assign v_RD_13590_out0 = v_RDN_4519_out0;
assign v_RD_13591_out0 = v_RDN_4520_out0;
assign v_RD_13592_out0 = v_RDN_4521_out0;
assign v_RD_13593_out0 = v_RDN_4522_out0;
assign v_RD_13594_out0 = v_RDN_4523_out0;
assign v_RD_13595_out0 = v_RDN_4524_out0;
assign v_RD_13596_out0 = v_RDN_4525_out0;
assign v_3_13619_out0 = v_B_3946_out0[3:3];
assign v_3_13620_out0 = v_B_3947_out0[3:3];
assign v_G14_13673_out0 = v_RD_13568_out0 && v__6831_out0;
assign v_G14_13674_out0 = v_RD_13569_out0 && v__6832_out0;
assign v_G14_13676_out0 = v_RD_13571_out0 && v__6834_out0;
assign v_G14_13688_out0 = v_RD_13583_out0 && v__6846_out0;
assign v_G14_13689_out0 = v_RD_13584_out0 && v__6847_out0;
assign v_G14_13691_out0 = v_RD_13586_out0 && v__6849_out0;
assign v__13770_out0 = { v_G7_8655_out0,v_G8_548_out0 };
assign v__13772_out0 = { v_G7_8657_out0,v_G8_550_out0 };
assign v__113_out0 = { v__386_out0,v__13770_out0 };
assign v__115_out0 = { v__388_out0,v__13772_out0 };
assign v_G15_132_out0 = v_RD_13567_out0 && v__1975_out0;
assign v_G15_135_out0 = v_RD_13570_out0 && v__1978_out0;
assign v_G15_137_out0 = v_RD_13572_out0 && v__1980_out0;
assign v_G15_138_out0 = v_RD_13573_out0 && v__1981_out0;
assign v_G15_139_out0 = v_RD_13574_out0 && v__1982_out0;
assign v_G15_140_out0 = v_RD_13575_out0 && v__1983_out0;
assign v_G15_141_out0 = v_RD_13576_out0 && v__1984_out0;
assign v_G15_142_out0 = v_RD_13577_out0 && v__1985_out0;
assign v_G15_143_out0 = v_RD_13578_out0 && v__1986_out0;
assign v_G15_144_out0 = v_RD_13579_out0 && v__1987_out0;
assign v_G15_145_out0 = v_RD_13580_out0 && v__1988_out0;
assign v_G15_146_out0 = v_RD_13581_out0 && v__1989_out0;
assign v_G15_147_out0 = v_RD_13582_out0 && v__1990_out0;
assign v_G15_150_out0 = v_RD_13585_out0 && v__1993_out0;
assign v_G15_152_out0 = v_RD_13587_out0 && v__1995_out0;
assign v_G15_153_out0 = v_RD_13588_out0 && v__1996_out0;
assign v_G15_154_out0 = v_RD_13589_out0 && v__1997_out0;
assign v_G15_155_out0 = v_RD_13590_out0 && v__1998_out0;
assign v_G15_156_out0 = v_RD_13591_out0 && v__1999_out0;
assign v_G15_157_out0 = v_RD_13592_out0 && v__2000_out0;
assign v_G15_158_out0 = v_RD_13593_out0 && v__2001_out0;
assign v_G15_159_out0 = v_RD_13594_out0 && v__2002_out0;
assign v_G15_160_out0 = v_RD_13595_out0 && v__2003_out0;
assign v_G15_161_out0 = v_RD_13596_out0 && v__2004_out0;
assign v__449_out0 = { v__7135_out0,v__2945_out0 };
assign v__451_out0 = { v__7137_out0,v__2947_out0 };
assign v_G5_638_out0 = ! v_EXP1_13488_out0;
assign v_G5_639_out0 = ! v_EXP1_13489_out0;
assign v_G11_651_out0 = v_RD_13567_out0 && v__3910_out0;
assign v_G11_654_out0 = v_RD_13570_out0 && v__3913_out0;
assign v_G11_656_out0 = v_RD_13572_out0 && v__3915_out0;
assign v_G11_657_out0 = v_RD_13573_out0 && v__3916_out0;
assign v_G11_658_out0 = v_RD_13574_out0 && v__3917_out0;
assign v_G11_659_out0 = v_RD_13575_out0 && v__3918_out0;
assign v_G11_660_out0 = v_RD_13576_out0 && v__3919_out0;
assign v_G11_661_out0 = v_RD_13577_out0 && v__3920_out0;
assign v_G11_662_out0 = v_RD_13578_out0 && v__3921_out0;
assign v_G11_663_out0 = v_RD_13579_out0 && v__3922_out0;
assign v_G11_664_out0 = v_RD_13580_out0 && v__3923_out0;
assign v_G11_665_out0 = v_RD_13581_out0 && v__3924_out0;
assign v_G11_666_out0 = v_RD_13582_out0 && v__3925_out0;
assign v_G11_669_out0 = v_RD_13585_out0 && v__3928_out0;
assign v_G11_671_out0 = v_RD_13587_out0 && v__3930_out0;
assign v_G11_672_out0 = v_RD_13588_out0 && v__3931_out0;
assign v_G11_673_out0 = v_RD_13589_out0 && v__3932_out0;
assign v_G11_674_out0 = v_RD_13590_out0 && v__3933_out0;
assign v_G11_675_out0 = v_RD_13591_out0 && v__3934_out0;
assign v_G11_676_out0 = v_RD_13592_out0 && v__3935_out0;
assign v_G11_677_out0 = v_RD_13593_out0 && v__3936_out0;
assign v_G11_678_out0 = v_RD_13594_out0 && v__3937_out0;
assign v_G11_679_out0 = v_RD_13595_out0 && v__3938_out0;
assign v_G11_680_out0 = v_RD_13596_out0 && v__3939_out0;
assign v__1212_out0 = { v__10456_out0,v_G16_11035_out0 };
assign v__1214_out0 = { v__10458_out0,v_G16_11037_out0 };
assign v__2345_out0 = { v__399_out0,v__13261_out0 };
assign v__2347_out0 = { v__401_out0,v__13263_out0 };
assign v__4733_out0 = { v__2649_out0,v_G11_2550_out0 };
assign v_RD_5874_out0 = v_G16_13183_out0;
assign v_RD_5897_out0 = v_RD_7204_out0;
assign v_RD_5899_out0 = v_RD_7205_out0;
assign v_RD_5904_out0 = v_G15_133_out0;
assign v_RD_5905_out0 = v_RD_7207_out0;
assign v_RD_5909_out0 = v_RD_7209_out0;
assign v_RD_5911_out0 = v_RD_7210_out0;
assign v_RD_5913_out0 = v_RD_7211_out0;
assign v_RD_5915_out0 = v_RD_7212_out0;
assign v_RD_5919_out0 = v_RD_7214_out0;
assign v_RD_5921_out0 = v_RD_7215_out0;
assign v_RD_5929_out0 = v_RD_7219_out0;
assign v_RD_5931_out0 = v_RD_7220_out0;
assign v_RD_5936_out0 = v_RD_7222_out0;
assign v_RD_5940_out0 = v_RD_7224_out0;
assign v_RD_5942_out0 = v_RD_7225_out0;
assign v_RD_5944_out0 = v_RD_7226_out0;
assign v_RD_5946_out0 = v_RD_7227_out0;
assign v_RD_5950_out0 = v_RD_7229_out0;
assign v_RD_5952_out0 = v_RD_7230_out0;
assign v_RD_5966_out0 = v_G16_13186_out0;
assign v_RD_5991_out0 = v_RD_7249_out0;
assign v_RD_5993_out0 = v_RD_7250_out0;
assign v_RD_5998_out0 = v_RD_7252_out0;
assign v_RD_6002_out0 = v_RD_7254_out0;
assign v_RD_6004_out0 = v_RD_7255_out0;
assign v_RD_6006_out0 = v_RD_7256_out0;
assign v_RD_6008_out0 = v_RD_7257_out0;
assign v_RD_6012_out0 = v_RD_7259_out0;
assign v_RD_6014_out0 = v_RD_7260_out0;
assign v_RD_6028_out0 = v_G16_13188_out0;
assign v_RD_6059_out0 = v_G16_13189_out0;
assign v_RD_6090_out0 = v_G16_13190_out0;
assign v_RD_6121_out0 = v_G16_13191_out0;
assign v_RD_6152_out0 = v_G16_13192_out0;
assign v_RD_6183_out0 = v_G16_13193_out0;
assign v_RD_6214_out0 = v_G16_13194_out0;
assign v_RD_6245_out0 = v_G16_13195_out0;
assign v_RD_6276_out0 = v_G16_13196_out0;
assign v_RD_6307_out0 = v_G16_13197_out0;
assign v_RD_6338_out0 = v_G16_13198_out0;
assign v_RD_6361_out0 = v_RD_7428_out0;
assign v_RD_6363_out0 = v_RD_7429_out0;
assign v_RD_6368_out0 = v_G15_148_out0;
assign v_RD_6369_out0 = v_RD_7431_out0;
assign v_RD_6373_out0 = v_RD_7433_out0;
assign v_RD_6375_out0 = v_RD_7434_out0;
assign v_RD_6377_out0 = v_RD_7435_out0;
assign v_RD_6379_out0 = v_RD_7436_out0;
assign v_RD_6383_out0 = v_RD_7438_out0;
assign v_RD_6385_out0 = v_RD_7439_out0;
assign v_RD_6393_out0 = v_RD_7443_out0;
assign v_RD_6395_out0 = v_RD_7444_out0;
assign v_RD_6400_out0 = v_RD_7446_out0;
assign v_RD_6404_out0 = v_RD_7448_out0;
assign v_RD_6406_out0 = v_RD_7449_out0;
assign v_RD_6408_out0 = v_RD_7450_out0;
assign v_RD_6410_out0 = v_RD_7451_out0;
assign v_RD_6414_out0 = v_RD_7453_out0;
assign v_RD_6416_out0 = v_RD_7454_out0;
assign v_RD_6430_out0 = v_G16_13201_out0;
assign v_RD_6455_out0 = v_RD_7473_out0;
assign v_RD_6457_out0 = v_RD_7474_out0;
assign v_RD_6462_out0 = v_RD_7476_out0;
assign v_RD_6466_out0 = v_RD_7478_out0;
assign v_RD_6468_out0 = v_RD_7479_out0;
assign v_RD_6470_out0 = v_RD_7480_out0;
assign v_RD_6472_out0 = v_RD_7481_out0;
assign v_RD_6476_out0 = v_RD_7483_out0;
assign v_RD_6478_out0 = v_RD_7484_out0;
assign v_RD_6492_out0 = v_G16_13203_out0;
assign v_RD_6523_out0 = v_G16_13204_out0;
assign v_RD_6554_out0 = v_G16_13205_out0;
assign v_RD_6585_out0 = v_G16_13206_out0;
assign v_RD_6616_out0 = v_G16_13207_out0;
assign v_RD_6647_out0 = v_G16_13208_out0;
assign v_RD_6678_out0 = v_G16_13209_out0;
assign v_RD_6709_out0 = v_G16_13210_out0;
assign v_RD_6740_out0 = v_G16_13211_out0;
assign v_RD_6771_out0 = v_G16_13212_out0;
assign v_G10_6975_out0 = v_RD_13567_out0 && v__2063_out0;
assign v_G10_6978_out0 = v_RD_13570_out0 && v__2066_out0;
assign v_G10_6980_out0 = v_RD_13572_out0 && v__2068_out0;
assign v_G10_6981_out0 = v_RD_13573_out0 && v__2069_out0;
assign v_G10_6982_out0 = v_RD_13574_out0 && v__2070_out0;
assign v_G10_6983_out0 = v_RD_13575_out0 && v__2071_out0;
assign v_G10_6984_out0 = v_RD_13576_out0 && v__2072_out0;
assign v_G10_6985_out0 = v_RD_13577_out0 && v__2073_out0;
assign v_G10_6986_out0 = v_RD_13578_out0 && v__2074_out0;
assign v_G10_6987_out0 = v_RD_13579_out0 && v__2075_out0;
assign v_G10_6988_out0 = v_RD_13580_out0 && v__2076_out0;
assign v_G10_6989_out0 = v_RD_13581_out0 && v__2077_out0;
assign v_G10_6990_out0 = v_RD_13582_out0 && v__2078_out0;
assign v_G10_6993_out0 = v_RD_13585_out0 && v__2081_out0;
assign v_G10_6995_out0 = v_RD_13587_out0 && v__2083_out0;
assign v_G10_6996_out0 = v_RD_13588_out0 && v__2084_out0;
assign v_G10_6997_out0 = v_RD_13589_out0 && v__2085_out0;
assign v_G10_6998_out0 = v_RD_13590_out0 && v__2086_out0;
assign v_G10_6999_out0 = v_RD_13591_out0 && v__2087_out0;
assign v_G10_7000_out0 = v_RD_13592_out0 && v__2088_out0;
assign v_G10_7001_out0 = v_RD_13593_out0 && v__2089_out0;
assign v_G10_7002_out0 = v_RD_13594_out0 && v__2090_out0;
assign v_G10_7003_out0 = v_RD_13595_out0 && v__2091_out0;
assign v_G10_7004_out0 = v_RD_13596_out0 && v__2092_out0;
assign v_RD_7190_out0 = v_G5_10621_out0;
assign v_RD_7191_out0 = v_G2_4620_out0;
assign v_RD_7193_out0 = v_G9_10572_out0;
assign v_RD_7195_out0 = v_G1_1909_out0;
assign v_RD_7196_out0 = v_G4_341_out0;
assign v_RD_7197_out0 = v_G6_2116_out0;
assign v_RD_7198_out0 = v_G7_11262_out0;
assign v_RD_7200_out0 = v_G8_2472_out0;
assign v_RD_7201_out0 = v_G3_241_out0;
assign v_RD_7202_out0 = v_G12_13222_out0;
assign v_RD_7203_out0 = v_G14_13673_out0;
assign v_RD_7206_out0 = v_G13_13353_out0;
assign v_RD_7208_out0 = v_G10_6976_out0;
assign v_RD_7213_out0 = v_G11_652_out0;
assign v_RD_7216_out0 = v_G12_13223_out0;
assign v_RD_7217_out0 = v_G14_13674_out0;
assign v_RD_7218_out0 = v_G15_134_out0;
assign v_RD_7221_out0 = v_G13_13354_out0;
assign v_RD_7223_out0 = v_G10_6977_out0;
assign v_RD_7228_out0 = v_G11_653_out0;
assign v_RD_7234_out0 = v_G5_10624_out0;
assign v_RD_7235_out0 = v_G2_4623_out0;
assign v_RD_7237_out0 = v_G9_10575_out0;
assign v_RD_7239_out0 = v_G1_1912_out0;
assign v_RD_7240_out0 = v_G4_344_out0;
assign v_RD_7241_out0 = v_G6_2119_out0;
assign v_RD_7242_out0 = v_G7_11265_out0;
assign v_RD_7244_out0 = v_G8_2475_out0;
assign v_RD_7245_out0 = v_G3_244_out0;
assign v_RD_7246_out0 = v_G12_13225_out0;
assign v_RD_7247_out0 = v_G14_13676_out0;
assign v_RD_7248_out0 = v_G15_136_out0;
assign v_RD_7251_out0 = v_G13_13356_out0;
assign v_RD_7253_out0 = v_G10_6979_out0;
assign v_RD_7258_out0 = v_G11_655_out0;
assign v_RD_7264_out0 = v_G5_10626_out0;
assign v_RD_7265_out0 = v_G2_4625_out0;
assign v_RD_7267_out0 = v_G9_10577_out0;
assign v_RD_7269_out0 = v_G1_1914_out0;
assign v_RD_7270_out0 = v_G4_346_out0;
assign v_RD_7271_out0 = v_G6_2121_out0;
assign v_RD_7272_out0 = v_G7_11267_out0;
assign v_RD_7274_out0 = v_G8_2477_out0;
assign v_RD_7275_out0 = v_G3_246_out0;
assign v_RD_7279_out0 = v_G5_10627_out0;
assign v_RD_7280_out0 = v_G2_4626_out0;
assign v_RD_7282_out0 = v_G9_10578_out0;
assign v_RD_7284_out0 = v_G1_1915_out0;
assign v_RD_7285_out0 = v_G4_347_out0;
assign v_RD_7286_out0 = v_G6_2122_out0;
assign v_RD_7287_out0 = v_G7_11268_out0;
assign v_RD_7289_out0 = v_G8_2478_out0;
assign v_RD_7290_out0 = v_G3_247_out0;
assign v_RD_7294_out0 = v_G5_10628_out0;
assign v_RD_7295_out0 = v_G2_4627_out0;
assign v_RD_7297_out0 = v_G9_10579_out0;
assign v_RD_7299_out0 = v_G1_1916_out0;
assign v_RD_7300_out0 = v_G4_348_out0;
assign v_RD_7301_out0 = v_G6_2123_out0;
assign v_RD_7302_out0 = v_G7_11269_out0;
assign v_RD_7304_out0 = v_G8_2479_out0;
assign v_RD_7305_out0 = v_G3_248_out0;
assign v_RD_7309_out0 = v_G5_10629_out0;
assign v_RD_7310_out0 = v_G2_4628_out0;
assign v_RD_7312_out0 = v_G9_10580_out0;
assign v_RD_7314_out0 = v_G1_1917_out0;
assign v_RD_7315_out0 = v_G4_349_out0;
assign v_RD_7316_out0 = v_G6_2124_out0;
assign v_RD_7317_out0 = v_G7_11270_out0;
assign v_RD_7319_out0 = v_G8_2480_out0;
assign v_RD_7320_out0 = v_G3_249_out0;
assign v_RD_7324_out0 = v_G5_10630_out0;
assign v_RD_7325_out0 = v_G2_4629_out0;
assign v_RD_7327_out0 = v_G9_10581_out0;
assign v_RD_7329_out0 = v_G1_1918_out0;
assign v_RD_7330_out0 = v_G4_350_out0;
assign v_RD_7331_out0 = v_G6_2125_out0;
assign v_RD_7332_out0 = v_G7_11271_out0;
assign v_RD_7334_out0 = v_G8_2481_out0;
assign v_RD_7335_out0 = v_G3_250_out0;
assign v_RD_7339_out0 = v_G5_10631_out0;
assign v_RD_7340_out0 = v_G2_4630_out0;
assign v_RD_7342_out0 = v_G9_10582_out0;
assign v_RD_7344_out0 = v_G1_1919_out0;
assign v_RD_7345_out0 = v_G4_351_out0;
assign v_RD_7346_out0 = v_G6_2126_out0;
assign v_RD_7347_out0 = v_G7_11272_out0;
assign v_RD_7349_out0 = v_G8_2482_out0;
assign v_RD_7350_out0 = v_G3_251_out0;
assign v_RD_7354_out0 = v_G5_10632_out0;
assign v_RD_7355_out0 = v_G2_4631_out0;
assign v_RD_7357_out0 = v_G9_10583_out0;
assign v_RD_7359_out0 = v_G1_1920_out0;
assign v_RD_7360_out0 = v_G4_352_out0;
assign v_RD_7361_out0 = v_G6_2127_out0;
assign v_RD_7362_out0 = v_G7_11273_out0;
assign v_RD_7364_out0 = v_G8_2483_out0;
assign v_RD_7365_out0 = v_G3_252_out0;
assign v_RD_7369_out0 = v_G5_10633_out0;
assign v_RD_7370_out0 = v_G2_4632_out0;
assign v_RD_7372_out0 = v_G9_10584_out0;
assign v_RD_7374_out0 = v_G1_1921_out0;
assign v_RD_7375_out0 = v_G4_353_out0;
assign v_RD_7376_out0 = v_G6_2128_out0;
assign v_RD_7377_out0 = v_G7_11274_out0;
assign v_RD_7379_out0 = v_G8_2484_out0;
assign v_RD_7380_out0 = v_G3_253_out0;
assign v_RD_7384_out0 = v_G5_10634_out0;
assign v_RD_7385_out0 = v_G2_4633_out0;
assign v_RD_7387_out0 = v_G9_10585_out0;
assign v_RD_7389_out0 = v_G1_1922_out0;
assign v_RD_7390_out0 = v_G4_354_out0;
assign v_RD_7391_out0 = v_G6_2129_out0;
assign v_RD_7392_out0 = v_G7_11275_out0;
assign v_RD_7394_out0 = v_G8_2485_out0;
assign v_RD_7395_out0 = v_G3_254_out0;
assign v_RD_7399_out0 = v_G5_10635_out0;
assign v_RD_7400_out0 = v_G2_4634_out0;
assign v_RD_7402_out0 = v_G9_10586_out0;
assign v_RD_7404_out0 = v_G1_1923_out0;
assign v_RD_7405_out0 = v_G4_355_out0;
assign v_RD_7406_out0 = v_G6_2130_out0;
assign v_RD_7407_out0 = v_G7_11276_out0;
assign v_RD_7409_out0 = v_G8_2486_out0;
assign v_RD_7410_out0 = v_G3_255_out0;
assign v_RD_7414_out0 = v_G5_10636_out0;
assign v_RD_7415_out0 = v_G2_4635_out0;
assign v_RD_7417_out0 = v_G9_10587_out0;
assign v_RD_7419_out0 = v_G1_1924_out0;
assign v_RD_7420_out0 = v_G4_356_out0;
assign v_RD_7421_out0 = v_G6_2131_out0;
assign v_RD_7422_out0 = v_G7_11277_out0;
assign v_RD_7424_out0 = v_G8_2487_out0;
assign v_RD_7425_out0 = v_G3_256_out0;
assign v_RD_7426_out0 = v_G12_13237_out0;
assign v_RD_7427_out0 = v_G14_13688_out0;
assign v_RD_7430_out0 = v_G13_13368_out0;
assign v_RD_7432_out0 = v_G10_6991_out0;
assign v_RD_7437_out0 = v_G11_667_out0;
assign v_RD_7440_out0 = v_G12_13238_out0;
assign v_RD_7441_out0 = v_G14_13689_out0;
assign v_RD_7442_out0 = v_G15_149_out0;
assign v_RD_7445_out0 = v_G13_13369_out0;
assign v_RD_7447_out0 = v_G10_6992_out0;
assign v_RD_7452_out0 = v_G11_668_out0;
assign v_RD_7458_out0 = v_G5_10639_out0;
assign v_RD_7459_out0 = v_G2_4638_out0;
assign v_RD_7461_out0 = v_G9_10590_out0;
assign v_RD_7463_out0 = v_G1_1927_out0;
assign v_RD_7464_out0 = v_G4_359_out0;
assign v_RD_7465_out0 = v_G6_2134_out0;
assign v_RD_7466_out0 = v_G7_11280_out0;
assign v_RD_7468_out0 = v_G8_2490_out0;
assign v_RD_7469_out0 = v_G3_259_out0;
assign v_RD_7470_out0 = v_G12_13240_out0;
assign v_RD_7471_out0 = v_G14_13691_out0;
assign v_RD_7472_out0 = v_G15_151_out0;
assign v_RD_7475_out0 = v_G13_13371_out0;
assign v_RD_7477_out0 = v_G10_6994_out0;
assign v_RD_7482_out0 = v_G11_670_out0;
assign v_RD_7488_out0 = v_G5_10641_out0;
assign v_RD_7489_out0 = v_G2_4640_out0;
assign v_RD_7491_out0 = v_G9_10592_out0;
assign v_RD_7493_out0 = v_G1_1929_out0;
assign v_RD_7494_out0 = v_G4_361_out0;
assign v_RD_7495_out0 = v_G6_2136_out0;
assign v_RD_7496_out0 = v_G7_11282_out0;
assign v_RD_7498_out0 = v_G8_2492_out0;
assign v_RD_7499_out0 = v_G3_261_out0;
assign v_RD_7503_out0 = v_G5_10642_out0;
assign v_RD_7504_out0 = v_G2_4641_out0;
assign v_RD_7506_out0 = v_G9_10593_out0;
assign v_RD_7508_out0 = v_G1_1930_out0;
assign v_RD_7509_out0 = v_G4_362_out0;
assign v_RD_7510_out0 = v_G6_2137_out0;
assign v_RD_7511_out0 = v_G7_11283_out0;
assign v_RD_7513_out0 = v_G8_2493_out0;
assign v_RD_7514_out0 = v_G3_262_out0;
assign v_RD_7518_out0 = v_G5_10643_out0;
assign v_RD_7519_out0 = v_G2_4642_out0;
assign v_RD_7521_out0 = v_G9_10594_out0;
assign v_RD_7523_out0 = v_G1_1931_out0;
assign v_RD_7524_out0 = v_G4_363_out0;
assign v_RD_7525_out0 = v_G6_2138_out0;
assign v_RD_7526_out0 = v_G7_11284_out0;
assign v_RD_7528_out0 = v_G8_2494_out0;
assign v_RD_7529_out0 = v_G3_263_out0;
assign v_RD_7533_out0 = v_G5_10644_out0;
assign v_RD_7534_out0 = v_G2_4643_out0;
assign v_RD_7536_out0 = v_G9_10595_out0;
assign v_RD_7538_out0 = v_G1_1932_out0;
assign v_RD_7539_out0 = v_G4_364_out0;
assign v_RD_7540_out0 = v_G6_2139_out0;
assign v_RD_7541_out0 = v_G7_11285_out0;
assign v_RD_7543_out0 = v_G8_2495_out0;
assign v_RD_7544_out0 = v_G3_264_out0;
assign v_RD_7548_out0 = v_G5_10645_out0;
assign v_RD_7549_out0 = v_G2_4644_out0;
assign v_RD_7551_out0 = v_G9_10596_out0;
assign v_RD_7553_out0 = v_G1_1933_out0;
assign v_RD_7554_out0 = v_G4_365_out0;
assign v_RD_7555_out0 = v_G6_2140_out0;
assign v_RD_7556_out0 = v_G7_11286_out0;
assign v_RD_7558_out0 = v_G8_2496_out0;
assign v_RD_7559_out0 = v_G3_265_out0;
assign v_RD_7563_out0 = v_G5_10646_out0;
assign v_RD_7564_out0 = v_G2_4645_out0;
assign v_RD_7566_out0 = v_G9_10597_out0;
assign v_RD_7568_out0 = v_G1_1934_out0;
assign v_RD_7569_out0 = v_G4_366_out0;
assign v_RD_7570_out0 = v_G6_2141_out0;
assign v_RD_7571_out0 = v_G7_11287_out0;
assign v_RD_7573_out0 = v_G8_2497_out0;
assign v_RD_7574_out0 = v_G3_266_out0;
assign v_RD_7578_out0 = v_G5_10647_out0;
assign v_RD_7579_out0 = v_G2_4646_out0;
assign v_RD_7581_out0 = v_G9_10598_out0;
assign v_RD_7583_out0 = v_G1_1935_out0;
assign v_RD_7584_out0 = v_G4_367_out0;
assign v_RD_7585_out0 = v_G6_2142_out0;
assign v_RD_7586_out0 = v_G7_11288_out0;
assign v_RD_7588_out0 = v_G8_2498_out0;
assign v_RD_7589_out0 = v_G3_267_out0;
assign v_RD_7593_out0 = v_G5_10648_out0;
assign v_RD_7594_out0 = v_G2_4647_out0;
assign v_RD_7596_out0 = v_G9_10599_out0;
assign v_RD_7598_out0 = v_G1_1936_out0;
assign v_RD_7599_out0 = v_G4_368_out0;
assign v_RD_7600_out0 = v_G6_2143_out0;
assign v_RD_7601_out0 = v_G7_11289_out0;
assign v_RD_7603_out0 = v_G8_2499_out0;
assign v_RD_7604_out0 = v_G3_268_out0;
assign v_RD_7608_out0 = v_G5_10649_out0;
assign v_RD_7609_out0 = v_G2_4648_out0;
assign v_RD_7611_out0 = v_G9_10600_out0;
assign v_RD_7613_out0 = v_G1_1937_out0;
assign v_RD_7614_out0 = v_G4_369_out0;
assign v_RD_7615_out0 = v_G6_2144_out0;
assign v_RD_7616_out0 = v_G7_11290_out0;
assign v_RD_7618_out0 = v_G8_2500_out0;
assign v_RD_7619_out0 = v_G3_269_out0;
assign v_RD_7623_out0 = v_G5_10650_out0;
assign v_RD_7624_out0 = v_G2_4649_out0;
assign v_RD_7626_out0 = v_G9_10601_out0;
assign v_RD_7628_out0 = v_G1_1938_out0;
assign v_RD_7629_out0 = v_G4_370_out0;
assign v_RD_7630_out0 = v_G6_2145_out0;
assign v_RD_7631_out0 = v_G7_11291_out0;
assign v_RD_7633_out0 = v_G8_2501_out0;
assign v_RD_7634_out0 = v_G3_270_out0;
assign v_IN_8838_out0 = v_IN_10403_out0;
assign v_IN_8839_out0 = v_IN_10404_out0;
assign v__10372_out0 = { v__3215_out0,v__3278_out0 };
assign v__10374_out0 = { v__3217_out0,v__3280_out0 };
assign v__11049_out0 = v_IN_10403_out0[13:0];
assign v__11049_out1 = v_IN_10403_out0[15:2];
assign v__11050_out0 = v_IN_10404_out0[13:0];
assign v__11050_out1 = v_IN_10404_out0[15:2];
assign v_G12_13221_out0 = v_RD_13567_out0 && v__2273_out0;
assign v_G12_13224_out0 = v_RD_13570_out0 && v__2276_out0;
assign v_G12_13226_out0 = v_RD_13572_out0 && v__2278_out0;
assign v_G12_13227_out0 = v_RD_13573_out0 && v__2279_out0;
assign v_G12_13228_out0 = v_RD_13574_out0 && v__2280_out0;
assign v_G12_13229_out0 = v_RD_13575_out0 && v__2281_out0;
assign v_G12_13230_out0 = v_RD_13576_out0 && v__2282_out0;
assign v_G12_13231_out0 = v_RD_13577_out0 && v__2283_out0;
assign v_G12_13232_out0 = v_RD_13578_out0 && v__2284_out0;
assign v_G12_13233_out0 = v_RD_13579_out0 && v__2285_out0;
assign v_G12_13234_out0 = v_RD_13580_out0 && v__2286_out0;
assign v_G12_13235_out0 = v_RD_13581_out0 && v__2287_out0;
assign v_G12_13236_out0 = v_RD_13582_out0 && v__2288_out0;
assign v_G12_13239_out0 = v_RD_13585_out0 && v__2291_out0;
assign v_G12_13241_out0 = v_RD_13587_out0 && v__2293_out0;
assign v_G12_13242_out0 = v_RD_13588_out0 && v__2294_out0;
assign v_G12_13243_out0 = v_RD_13589_out0 && v__2295_out0;
assign v_G12_13244_out0 = v_RD_13590_out0 && v__2296_out0;
assign v_G12_13245_out0 = v_RD_13591_out0 && v__2297_out0;
assign v_G12_13246_out0 = v_RD_13592_out0 && v__2298_out0;
assign v_G12_13247_out0 = v_RD_13593_out0 && v__2299_out0;
assign v_G12_13248_out0 = v_RD_13594_out0 && v__2300_out0;
assign v_G12_13249_out0 = v_RD_13595_out0 && v__2301_out0;
assign v_G12_13250_out0 = v_RD_13596_out0 && v__2302_out0;
assign v_G13_13352_out0 = v_RD_13567_out0 && v__13715_out0;
assign v_G13_13355_out0 = v_RD_13570_out0 && v__13718_out0;
assign v_G13_13357_out0 = v_RD_13572_out0 && v__13720_out0;
assign v_G13_13358_out0 = v_RD_13573_out0 && v__13721_out0;
assign v_G13_13359_out0 = v_RD_13574_out0 && v__13722_out0;
assign v_G13_13360_out0 = v_RD_13575_out0 && v__13723_out0;
assign v_G13_13361_out0 = v_RD_13576_out0 && v__13724_out0;
assign v_G13_13362_out0 = v_RD_13577_out0 && v__13725_out0;
assign v_G13_13363_out0 = v_RD_13578_out0 && v__13726_out0;
assign v_G13_13364_out0 = v_RD_13579_out0 && v__13727_out0;
assign v_G13_13365_out0 = v_RD_13580_out0 && v__13728_out0;
assign v_G13_13366_out0 = v_RD_13581_out0 && v__13729_out0;
assign v_G13_13367_out0 = v_RD_13582_out0 && v__13730_out0;
assign v_G13_13370_out0 = v_RD_13585_out0 && v__13733_out0;
assign v_G13_13372_out0 = v_RD_13587_out0 && v__13735_out0;
assign v_G13_13373_out0 = v_RD_13588_out0 && v__13736_out0;
assign v_G13_13374_out0 = v_RD_13589_out0 && v__13737_out0;
assign v_G13_13375_out0 = v_RD_13590_out0 && v__13738_out0;
assign v_G13_13376_out0 = v_RD_13591_out0 && v__13739_out0;
assign v_G13_13377_out0 = v_RD_13592_out0 && v__13740_out0;
assign v_G13_13378_out0 = v_RD_13593_out0 && v__13741_out0;
assign v_G13_13379_out0 = v_RD_13594_out0 && v__13742_out0;
assign v_G13_13380_out0 = v_RD_13595_out0 && v__13743_out0;
assign v_G13_13381_out0 = v_RD_13596_out0 && v__13744_out0;
assign v_IN_13668_out0 = v_SIG_TO_SHIFT_5836_out0;
assign v_IN_13669_out0 = v_SIG_TO_SHIFT_5837_out0;
assign v_G14_13672_out0 = v_RD_13567_out0 && v__6830_out0;
assign v_G14_13675_out0 = v_RD_13570_out0 && v__6833_out0;
assign v_G14_13677_out0 = v_RD_13572_out0 && v__6835_out0;
assign v_G14_13678_out0 = v_RD_13573_out0 && v__6836_out0;
assign v_G14_13679_out0 = v_RD_13574_out0 && v__6837_out0;
assign v_G14_13680_out0 = v_RD_13575_out0 && v__6838_out0;
assign v_G14_13681_out0 = v_RD_13576_out0 && v__6839_out0;
assign v_G14_13682_out0 = v_RD_13577_out0 && v__6840_out0;
assign v_G14_13683_out0 = v_RD_13578_out0 && v__6841_out0;
assign v_G14_13684_out0 = v_RD_13579_out0 && v__6842_out0;
assign v_G14_13685_out0 = v_RD_13580_out0 && v__6843_out0;
assign v_G14_13686_out0 = v_RD_13581_out0 && v__6844_out0;
assign v_G14_13687_out0 = v_RD_13582_out0 && v__6845_out0;
assign v_G14_13690_out0 = v_RD_13585_out0 && v__6848_out0;
assign v_G14_13692_out0 = v_RD_13587_out0 && v__6850_out0;
assign v_G14_13693_out0 = v_RD_13588_out0 && v__6851_out0;
assign v_G14_13694_out0 = v_RD_13589_out0 && v__6852_out0;
assign v_G14_13695_out0 = v_RD_13590_out0 && v__6853_out0;
assign v_G14_13696_out0 = v_RD_13591_out0 && v__6854_out0;
assign v_G14_13697_out0 = v_RD_13592_out0 && v__6855_out0;
assign v_G14_13698_out0 = v_RD_13593_out0 && v__6856_out0;
assign v_G14_13699_out0 = v_RD_13594_out0 && v__6857_out0;
assign v_G14_13700_out0 = v_RD_13595_out0 && v__6858_out0;
assign v_G14_13701_out0 = v_RD_13596_out0 && v__6859_out0;
assign v_IN1_2189_out0 = v_IN_13668_out0;
assign v_IN1_2190_out0 = v_IN_13669_out0;
assign v_NOTUSED_2589_out0 = v__11049_out1;
assign v_NOTUSED_2590_out0 = v__11050_out1;
assign v__2684_out0 = { v__10372_out0,v__113_out0 };
assign v__2686_out0 = { v__10374_out0,v__115_out0 };
assign v__4449_out0 = { v__2345_out0,v__449_out0 };
assign v__4451_out0 = { v__2347_out0,v__451_out0 };
assign v_RD_5868_out0 = v_RD_7190_out0;
assign v_RD_5870_out0 = v_RD_7191_out0;
assign v_RD_5875_out0 = v_RD_7193_out0;
assign v_RD_5879_out0 = v_RD_7195_out0;
assign v_RD_5881_out0 = v_RD_7196_out0;
assign v_RD_5883_out0 = v_RD_7197_out0;
assign v_RD_5885_out0 = v_RD_7198_out0;
assign v_RD_5889_out0 = v_RD_7200_out0;
assign v_RD_5891_out0 = v_RD_7201_out0;
assign v_RD_5893_out0 = v_RD_7202_out0;
assign v_RD_5895_out0 = v_RD_7203_out0;
assign v_RD_5901_out0 = v_RD_7206_out0;
assign v_RD_5907_out0 = v_RD_7208_out0;
assign v_RD_5917_out0 = v_RD_7213_out0;
assign v_RD_5923_out0 = v_RD_7216_out0;
assign v_RD_5925_out0 = v_RD_7217_out0;
assign v_RD_5927_out0 = v_RD_7218_out0;
assign v_RD_5933_out0 = v_RD_7221_out0;
assign v_RD_5938_out0 = v_RD_7223_out0;
assign v_RD_5948_out0 = v_RD_7228_out0;
assign v_RD_5960_out0 = v_RD_7234_out0;
assign v_RD_5962_out0 = v_RD_7235_out0;
assign v_RD_5967_out0 = v_RD_7237_out0;
assign v_RD_5971_out0 = v_RD_7239_out0;
assign v_RD_5973_out0 = v_RD_7240_out0;
assign v_RD_5975_out0 = v_RD_7241_out0;
assign v_RD_5977_out0 = v_RD_7242_out0;
assign v_RD_5981_out0 = v_RD_7244_out0;
assign v_RD_5983_out0 = v_RD_7245_out0;
assign v_RD_5985_out0 = v_RD_7246_out0;
assign v_RD_5987_out0 = v_RD_7247_out0;
assign v_RD_5989_out0 = v_RD_7248_out0;
assign v_RD_5995_out0 = v_RD_7251_out0;
assign v_RD_6000_out0 = v_RD_7253_out0;
assign v_RD_6010_out0 = v_RD_7258_out0;
assign v_RD_6022_out0 = v_RD_7264_out0;
assign v_RD_6024_out0 = v_RD_7265_out0;
assign v_RD_6029_out0 = v_RD_7267_out0;
assign v_RD_6033_out0 = v_RD_7269_out0;
assign v_RD_6035_out0 = v_RD_7270_out0;
assign v_RD_6037_out0 = v_RD_7271_out0;
assign v_RD_6039_out0 = v_RD_7272_out0;
assign v_RD_6043_out0 = v_RD_7274_out0;
assign v_RD_6045_out0 = v_RD_7275_out0;
assign v_RD_6053_out0 = v_RD_7279_out0;
assign v_RD_6055_out0 = v_RD_7280_out0;
assign v_RD_6060_out0 = v_RD_7282_out0;
assign v_RD_6064_out0 = v_RD_7284_out0;
assign v_RD_6066_out0 = v_RD_7285_out0;
assign v_RD_6068_out0 = v_RD_7286_out0;
assign v_RD_6070_out0 = v_RD_7287_out0;
assign v_RD_6074_out0 = v_RD_7289_out0;
assign v_RD_6076_out0 = v_RD_7290_out0;
assign v_RD_6084_out0 = v_RD_7294_out0;
assign v_RD_6086_out0 = v_RD_7295_out0;
assign v_RD_6091_out0 = v_RD_7297_out0;
assign v_RD_6095_out0 = v_RD_7299_out0;
assign v_RD_6097_out0 = v_RD_7300_out0;
assign v_RD_6099_out0 = v_RD_7301_out0;
assign v_RD_6101_out0 = v_RD_7302_out0;
assign v_RD_6105_out0 = v_RD_7304_out0;
assign v_RD_6107_out0 = v_RD_7305_out0;
assign v_RD_6115_out0 = v_RD_7309_out0;
assign v_RD_6117_out0 = v_RD_7310_out0;
assign v_RD_6122_out0 = v_RD_7312_out0;
assign v_RD_6126_out0 = v_RD_7314_out0;
assign v_RD_6128_out0 = v_RD_7315_out0;
assign v_RD_6130_out0 = v_RD_7316_out0;
assign v_RD_6132_out0 = v_RD_7317_out0;
assign v_RD_6136_out0 = v_RD_7319_out0;
assign v_RD_6138_out0 = v_RD_7320_out0;
assign v_RD_6146_out0 = v_RD_7324_out0;
assign v_RD_6148_out0 = v_RD_7325_out0;
assign v_RD_6153_out0 = v_RD_7327_out0;
assign v_RD_6157_out0 = v_RD_7329_out0;
assign v_RD_6159_out0 = v_RD_7330_out0;
assign v_RD_6161_out0 = v_RD_7331_out0;
assign v_RD_6163_out0 = v_RD_7332_out0;
assign v_RD_6167_out0 = v_RD_7334_out0;
assign v_RD_6169_out0 = v_RD_7335_out0;
assign v_RD_6177_out0 = v_RD_7339_out0;
assign v_RD_6179_out0 = v_RD_7340_out0;
assign v_RD_6184_out0 = v_RD_7342_out0;
assign v_RD_6188_out0 = v_RD_7344_out0;
assign v_RD_6190_out0 = v_RD_7345_out0;
assign v_RD_6192_out0 = v_RD_7346_out0;
assign v_RD_6194_out0 = v_RD_7347_out0;
assign v_RD_6198_out0 = v_RD_7349_out0;
assign v_RD_6200_out0 = v_RD_7350_out0;
assign v_RD_6208_out0 = v_RD_7354_out0;
assign v_RD_6210_out0 = v_RD_7355_out0;
assign v_RD_6215_out0 = v_RD_7357_out0;
assign v_RD_6219_out0 = v_RD_7359_out0;
assign v_RD_6221_out0 = v_RD_7360_out0;
assign v_RD_6223_out0 = v_RD_7361_out0;
assign v_RD_6225_out0 = v_RD_7362_out0;
assign v_RD_6229_out0 = v_RD_7364_out0;
assign v_RD_6231_out0 = v_RD_7365_out0;
assign v_RD_6239_out0 = v_RD_7369_out0;
assign v_RD_6241_out0 = v_RD_7370_out0;
assign v_RD_6246_out0 = v_RD_7372_out0;
assign v_RD_6250_out0 = v_RD_7374_out0;
assign v_RD_6252_out0 = v_RD_7375_out0;
assign v_RD_6254_out0 = v_RD_7376_out0;
assign v_RD_6256_out0 = v_RD_7377_out0;
assign v_RD_6260_out0 = v_RD_7379_out0;
assign v_RD_6262_out0 = v_RD_7380_out0;
assign v_RD_6270_out0 = v_RD_7384_out0;
assign v_RD_6272_out0 = v_RD_7385_out0;
assign v_RD_6277_out0 = v_RD_7387_out0;
assign v_RD_6281_out0 = v_RD_7389_out0;
assign v_RD_6283_out0 = v_RD_7390_out0;
assign v_RD_6285_out0 = v_RD_7391_out0;
assign v_RD_6287_out0 = v_RD_7392_out0;
assign v_RD_6291_out0 = v_RD_7394_out0;
assign v_RD_6293_out0 = v_RD_7395_out0;
assign v_RD_6301_out0 = v_RD_7399_out0;
assign v_RD_6303_out0 = v_RD_7400_out0;
assign v_RD_6308_out0 = v_RD_7402_out0;
assign v_RD_6312_out0 = v_RD_7404_out0;
assign v_RD_6314_out0 = v_RD_7405_out0;
assign v_RD_6316_out0 = v_RD_7406_out0;
assign v_RD_6318_out0 = v_RD_7407_out0;
assign v_RD_6322_out0 = v_RD_7409_out0;
assign v_RD_6324_out0 = v_RD_7410_out0;
assign v_RD_6332_out0 = v_RD_7414_out0;
assign v_RD_6334_out0 = v_RD_7415_out0;
assign v_RD_6339_out0 = v_RD_7417_out0;
assign v_RD_6343_out0 = v_RD_7419_out0;
assign v_RD_6345_out0 = v_RD_7420_out0;
assign v_RD_6347_out0 = v_RD_7421_out0;
assign v_RD_6349_out0 = v_RD_7422_out0;
assign v_RD_6353_out0 = v_RD_7424_out0;
assign v_RD_6355_out0 = v_RD_7425_out0;
assign v_RD_6357_out0 = v_RD_7426_out0;
assign v_RD_6359_out0 = v_RD_7427_out0;
assign v_RD_6365_out0 = v_RD_7430_out0;
assign v_RD_6371_out0 = v_RD_7432_out0;
assign v_RD_6381_out0 = v_RD_7437_out0;
assign v_RD_6387_out0 = v_RD_7440_out0;
assign v_RD_6389_out0 = v_RD_7441_out0;
assign v_RD_6391_out0 = v_RD_7442_out0;
assign v_RD_6397_out0 = v_RD_7445_out0;
assign v_RD_6402_out0 = v_RD_7447_out0;
assign v_RD_6412_out0 = v_RD_7452_out0;
assign v_RD_6424_out0 = v_RD_7458_out0;
assign v_RD_6426_out0 = v_RD_7459_out0;
assign v_RD_6431_out0 = v_RD_7461_out0;
assign v_RD_6435_out0 = v_RD_7463_out0;
assign v_RD_6437_out0 = v_RD_7464_out0;
assign v_RD_6439_out0 = v_RD_7465_out0;
assign v_RD_6441_out0 = v_RD_7466_out0;
assign v_RD_6445_out0 = v_RD_7468_out0;
assign v_RD_6447_out0 = v_RD_7469_out0;
assign v_RD_6449_out0 = v_RD_7470_out0;
assign v_RD_6451_out0 = v_RD_7471_out0;
assign v_RD_6453_out0 = v_RD_7472_out0;
assign v_RD_6459_out0 = v_RD_7475_out0;
assign v_RD_6464_out0 = v_RD_7477_out0;
assign v_RD_6474_out0 = v_RD_7482_out0;
assign v_RD_6486_out0 = v_RD_7488_out0;
assign v_RD_6488_out0 = v_RD_7489_out0;
assign v_RD_6493_out0 = v_RD_7491_out0;
assign v_RD_6497_out0 = v_RD_7493_out0;
assign v_RD_6499_out0 = v_RD_7494_out0;
assign v_RD_6501_out0 = v_RD_7495_out0;
assign v_RD_6503_out0 = v_RD_7496_out0;
assign v_RD_6507_out0 = v_RD_7498_out0;
assign v_RD_6509_out0 = v_RD_7499_out0;
assign v_RD_6517_out0 = v_RD_7503_out0;
assign v_RD_6519_out0 = v_RD_7504_out0;
assign v_RD_6524_out0 = v_RD_7506_out0;
assign v_RD_6528_out0 = v_RD_7508_out0;
assign v_RD_6530_out0 = v_RD_7509_out0;
assign v_RD_6532_out0 = v_RD_7510_out0;
assign v_RD_6534_out0 = v_RD_7511_out0;
assign v_RD_6538_out0 = v_RD_7513_out0;
assign v_RD_6540_out0 = v_RD_7514_out0;
assign v_RD_6548_out0 = v_RD_7518_out0;
assign v_RD_6550_out0 = v_RD_7519_out0;
assign v_RD_6555_out0 = v_RD_7521_out0;
assign v_RD_6559_out0 = v_RD_7523_out0;
assign v_RD_6561_out0 = v_RD_7524_out0;
assign v_RD_6563_out0 = v_RD_7525_out0;
assign v_RD_6565_out0 = v_RD_7526_out0;
assign v_RD_6569_out0 = v_RD_7528_out0;
assign v_RD_6571_out0 = v_RD_7529_out0;
assign v_RD_6579_out0 = v_RD_7533_out0;
assign v_RD_6581_out0 = v_RD_7534_out0;
assign v_RD_6586_out0 = v_RD_7536_out0;
assign v_RD_6590_out0 = v_RD_7538_out0;
assign v_RD_6592_out0 = v_RD_7539_out0;
assign v_RD_6594_out0 = v_RD_7540_out0;
assign v_RD_6596_out0 = v_RD_7541_out0;
assign v_RD_6600_out0 = v_RD_7543_out0;
assign v_RD_6602_out0 = v_RD_7544_out0;
assign v_RD_6610_out0 = v_RD_7548_out0;
assign v_RD_6612_out0 = v_RD_7549_out0;
assign v_RD_6617_out0 = v_RD_7551_out0;
assign v_RD_6621_out0 = v_RD_7553_out0;
assign v_RD_6623_out0 = v_RD_7554_out0;
assign v_RD_6625_out0 = v_RD_7555_out0;
assign v_RD_6627_out0 = v_RD_7556_out0;
assign v_RD_6631_out0 = v_RD_7558_out0;
assign v_RD_6633_out0 = v_RD_7559_out0;
assign v_RD_6641_out0 = v_RD_7563_out0;
assign v_RD_6643_out0 = v_RD_7564_out0;
assign v_RD_6648_out0 = v_RD_7566_out0;
assign v_RD_6652_out0 = v_RD_7568_out0;
assign v_RD_6654_out0 = v_RD_7569_out0;
assign v_RD_6656_out0 = v_RD_7570_out0;
assign v_RD_6658_out0 = v_RD_7571_out0;
assign v_RD_6662_out0 = v_RD_7573_out0;
assign v_RD_6664_out0 = v_RD_7574_out0;
assign v_RD_6672_out0 = v_RD_7578_out0;
assign v_RD_6674_out0 = v_RD_7579_out0;
assign v_RD_6679_out0 = v_RD_7581_out0;
assign v_RD_6683_out0 = v_RD_7583_out0;
assign v_RD_6685_out0 = v_RD_7584_out0;
assign v_RD_6687_out0 = v_RD_7585_out0;
assign v_RD_6689_out0 = v_RD_7586_out0;
assign v_RD_6693_out0 = v_RD_7588_out0;
assign v_RD_6695_out0 = v_RD_7589_out0;
assign v_RD_6703_out0 = v_RD_7593_out0;
assign v_RD_6705_out0 = v_RD_7594_out0;
assign v_RD_6710_out0 = v_RD_7596_out0;
assign v_RD_6714_out0 = v_RD_7598_out0;
assign v_RD_6716_out0 = v_RD_7599_out0;
assign v_RD_6718_out0 = v_RD_7600_out0;
assign v_RD_6720_out0 = v_RD_7601_out0;
assign v_RD_6724_out0 = v_RD_7603_out0;
assign v_RD_6726_out0 = v_RD_7604_out0;
assign v_RD_6734_out0 = v_RD_7608_out0;
assign v_RD_6736_out0 = v_RD_7609_out0;
assign v_RD_6741_out0 = v_RD_7611_out0;
assign v_RD_6745_out0 = v_RD_7613_out0;
assign v_RD_6747_out0 = v_RD_7614_out0;
assign v_RD_6749_out0 = v_RD_7615_out0;
assign v_RD_6751_out0 = v_RD_7616_out0;
assign v_RD_6755_out0 = v_RD_7618_out0;
assign v_RD_6757_out0 = v_RD_7619_out0;
assign v_RD_6765_out0 = v_RD_7623_out0;
assign v_RD_6767_out0 = v_RD_7624_out0;
assign v_RD_6772_out0 = v_RD_7626_out0;
assign v_RD_6776_out0 = v_RD_7628_out0;
assign v_RD_6778_out0 = v_RD_7629_out0;
assign v_RD_6780_out0 = v_RD_7630_out0;
assign v_RD_6782_out0 = v_RD_7631_out0;
assign v_RD_6786_out0 = v_RD_7633_out0;
assign v_RD_6788_out0 = v_RD_7634_out0;
assign v_RD_7187_out0 = v_G12_13221_out0;
assign v_RD_7188_out0 = v_G14_13672_out0;
assign v_RD_7189_out0 = v_G15_132_out0;
assign v_RD_7192_out0 = v_G13_13352_out0;
assign v_RD_7194_out0 = v_G10_6975_out0;
assign v_RD_7199_out0 = v_G11_651_out0;
assign v_RD_7231_out0 = v_G12_13224_out0;
assign v_RD_7232_out0 = v_G14_13675_out0;
assign v_RD_7233_out0 = v_G15_135_out0;
assign v_RD_7236_out0 = v_G13_13355_out0;
assign v_RD_7238_out0 = v_G10_6978_out0;
assign v_RD_7243_out0 = v_G11_654_out0;
assign v_RD_7261_out0 = v_G12_13226_out0;
assign v_RD_7262_out0 = v_G14_13677_out0;
assign v_RD_7263_out0 = v_G15_137_out0;
assign v_RD_7266_out0 = v_G13_13357_out0;
assign v_RD_7268_out0 = v_G10_6980_out0;
assign v_RD_7273_out0 = v_G11_656_out0;
assign v_RD_7276_out0 = v_G12_13227_out0;
assign v_RD_7277_out0 = v_G14_13678_out0;
assign v_RD_7278_out0 = v_G15_138_out0;
assign v_RD_7281_out0 = v_G13_13358_out0;
assign v_RD_7283_out0 = v_G10_6981_out0;
assign v_RD_7288_out0 = v_G11_657_out0;
assign v_RD_7291_out0 = v_G12_13228_out0;
assign v_RD_7292_out0 = v_G14_13679_out0;
assign v_RD_7293_out0 = v_G15_139_out0;
assign v_RD_7296_out0 = v_G13_13359_out0;
assign v_RD_7298_out0 = v_G10_6982_out0;
assign v_RD_7303_out0 = v_G11_658_out0;
assign v_RD_7306_out0 = v_G12_13229_out0;
assign v_RD_7307_out0 = v_G14_13680_out0;
assign v_RD_7308_out0 = v_G15_140_out0;
assign v_RD_7311_out0 = v_G13_13360_out0;
assign v_RD_7313_out0 = v_G10_6983_out0;
assign v_RD_7318_out0 = v_G11_659_out0;
assign v_RD_7321_out0 = v_G12_13230_out0;
assign v_RD_7322_out0 = v_G14_13681_out0;
assign v_RD_7323_out0 = v_G15_141_out0;
assign v_RD_7326_out0 = v_G13_13361_out0;
assign v_RD_7328_out0 = v_G10_6984_out0;
assign v_RD_7333_out0 = v_G11_660_out0;
assign v_RD_7336_out0 = v_G12_13231_out0;
assign v_RD_7337_out0 = v_G14_13682_out0;
assign v_RD_7338_out0 = v_G15_142_out0;
assign v_RD_7341_out0 = v_G13_13362_out0;
assign v_RD_7343_out0 = v_G10_6985_out0;
assign v_RD_7348_out0 = v_G11_661_out0;
assign v_RD_7351_out0 = v_G12_13232_out0;
assign v_RD_7352_out0 = v_G14_13683_out0;
assign v_RD_7353_out0 = v_G15_143_out0;
assign v_RD_7356_out0 = v_G13_13363_out0;
assign v_RD_7358_out0 = v_G10_6986_out0;
assign v_RD_7363_out0 = v_G11_662_out0;
assign v_RD_7366_out0 = v_G12_13233_out0;
assign v_RD_7367_out0 = v_G14_13684_out0;
assign v_RD_7368_out0 = v_G15_144_out0;
assign v_RD_7371_out0 = v_G13_13364_out0;
assign v_RD_7373_out0 = v_G10_6987_out0;
assign v_RD_7378_out0 = v_G11_663_out0;
assign v_RD_7381_out0 = v_G12_13234_out0;
assign v_RD_7382_out0 = v_G14_13685_out0;
assign v_RD_7383_out0 = v_G15_145_out0;
assign v_RD_7386_out0 = v_G13_13365_out0;
assign v_RD_7388_out0 = v_G10_6988_out0;
assign v_RD_7393_out0 = v_G11_664_out0;
assign v_RD_7396_out0 = v_G12_13235_out0;
assign v_RD_7397_out0 = v_G14_13686_out0;
assign v_RD_7398_out0 = v_G15_146_out0;
assign v_RD_7401_out0 = v_G13_13366_out0;
assign v_RD_7403_out0 = v_G10_6989_out0;
assign v_RD_7408_out0 = v_G11_665_out0;
assign v_RD_7411_out0 = v_G12_13236_out0;
assign v_RD_7412_out0 = v_G14_13687_out0;
assign v_RD_7413_out0 = v_G15_147_out0;
assign v_RD_7416_out0 = v_G13_13367_out0;
assign v_RD_7418_out0 = v_G10_6990_out0;
assign v_RD_7423_out0 = v_G11_666_out0;
assign v_RD_7455_out0 = v_G12_13239_out0;
assign v_RD_7456_out0 = v_G14_13690_out0;
assign v_RD_7457_out0 = v_G15_150_out0;
assign v_RD_7460_out0 = v_G13_13370_out0;
assign v_RD_7462_out0 = v_G10_6993_out0;
assign v_RD_7467_out0 = v_G11_669_out0;
assign v_RD_7485_out0 = v_G12_13241_out0;
assign v_RD_7486_out0 = v_G14_13692_out0;
assign v_RD_7487_out0 = v_G15_152_out0;
assign v_RD_7490_out0 = v_G13_13372_out0;
assign v_RD_7492_out0 = v_G10_6995_out0;
assign v_RD_7497_out0 = v_G11_671_out0;
assign v_RD_7500_out0 = v_G12_13242_out0;
assign v_RD_7501_out0 = v_G14_13693_out0;
assign v_RD_7502_out0 = v_G15_153_out0;
assign v_RD_7505_out0 = v_G13_13373_out0;
assign v_RD_7507_out0 = v_G10_6996_out0;
assign v_RD_7512_out0 = v_G11_672_out0;
assign v_RD_7515_out0 = v_G12_13243_out0;
assign v_RD_7516_out0 = v_G14_13694_out0;
assign v_RD_7517_out0 = v_G15_154_out0;
assign v_RD_7520_out0 = v_G13_13374_out0;
assign v_RD_7522_out0 = v_G10_6997_out0;
assign v_RD_7527_out0 = v_G11_673_out0;
assign v_RD_7530_out0 = v_G12_13244_out0;
assign v_RD_7531_out0 = v_G14_13695_out0;
assign v_RD_7532_out0 = v_G15_155_out0;
assign v_RD_7535_out0 = v_G13_13375_out0;
assign v_RD_7537_out0 = v_G10_6998_out0;
assign v_RD_7542_out0 = v_G11_674_out0;
assign v_RD_7545_out0 = v_G12_13245_out0;
assign v_RD_7546_out0 = v_G14_13696_out0;
assign v_RD_7547_out0 = v_G15_156_out0;
assign v_RD_7550_out0 = v_G13_13376_out0;
assign v_RD_7552_out0 = v_G10_6999_out0;
assign v_RD_7557_out0 = v_G11_675_out0;
assign v_RD_7560_out0 = v_G12_13246_out0;
assign v_RD_7561_out0 = v_G14_13697_out0;
assign v_RD_7562_out0 = v_G15_157_out0;
assign v_RD_7565_out0 = v_G13_13377_out0;
assign v_RD_7567_out0 = v_G10_7000_out0;
assign v_RD_7572_out0 = v_G11_676_out0;
assign v_RD_7575_out0 = v_G12_13247_out0;
assign v_RD_7576_out0 = v_G14_13698_out0;
assign v_RD_7577_out0 = v_G15_158_out0;
assign v_RD_7580_out0 = v_G13_13378_out0;
assign v_RD_7582_out0 = v_G10_7001_out0;
assign v_RD_7587_out0 = v_G11_677_out0;
assign v_RD_7590_out0 = v_G12_13248_out0;
assign v_RD_7591_out0 = v_G14_13699_out0;
assign v_RD_7592_out0 = v_G15_159_out0;
assign v_RD_7595_out0 = v_G13_13379_out0;
assign v_RD_7597_out0 = v_G10_7002_out0;
assign v_RD_7602_out0 = v_G11_678_out0;
assign v_RD_7605_out0 = v_G12_13249_out0;
assign v_RD_7606_out0 = v_G14_13700_out0;
assign v_RD_7607_out0 = v_G15_160_out0;
assign v_RD_7610_out0 = v_G13_13380_out0;
assign v_RD_7612_out0 = v_G10_7003_out0;
assign v_RD_7617_out0 = v_G11_679_out0;
assign v_RD_7620_out0 = v_G12_13250_out0;
assign v_RD_7621_out0 = v_G14_13701_out0;
assign v_RD_7622_out0 = v_G15_161_out0;
assign v_RD_7625_out0 = v_G13_13381_out0;
assign v_RD_7627_out0 = v_G10_7004_out0;
assign v_RD_7632_out0 = v_G11_680_out0;
assign v_ADDER_IN_8745_out0 = v__1212_out0;
assign v_ADDER_IN_8747_out0 = v__1214_out0;
assign v__10333_out0 = { v_C1_11292_out0,v__11049_out0 };
assign v__10334_out0 = { v_C1_11293_out0,v__11050_out0 };
assign v__10783_out0 = { v__4733_out0,v_G12_4699_out0 };
assign v_MUX1_6_out0 = v_LSL_2842_out0 ? v__10333_out0 : v_IN_8838_out0;
assign v_MUX1_7_out0 = v_LSL_2843_out0 ? v__10334_out0 : v_IN_8839_out0;
assign v__1867_out0 = { v__2684_out0,v__4449_out0 };
assign v__1869_out0 = { v__2686_out0,v__4451_out0 };
assign {v_A1_3174_out1,v_A1_3174_out0 } = v_RM_13508_out0 + v_ADDER_IN_8745_out0 + v_U_10469_out0;
assign {v_A1_3175_out1,v_A1_3175_out0 } = v_RM_13509_out0 + v_ADDER_IN_8747_out0 + v_U_10470_out0;
assign v__3907_out0 = v_IN1_2189_out0[0:0];
assign v__3907_out1 = v_IN1_2189_out0[10:10];
assign v__3908_out0 = v_IN1_2190_out0[0:0];
assign v__3908_out1 = v_IN1_2190_out0[10:10];
assign v_RD_5862_out0 = v_RD_7187_out0;
assign v_RD_5864_out0 = v_RD_7188_out0;
assign v_RD_5866_out0 = v_RD_7189_out0;
assign v_RD_5872_out0 = v_RD_7192_out0;
assign v_RD_5877_out0 = v_RD_7194_out0;
assign v_RD_5887_out0 = v_RD_7199_out0;
assign v_RD_5954_out0 = v_RD_7231_out0;
assign v_RD_5956_out0 = v_RD_7232_out0;
assign v_RD_5958_out0 = v_RD_7233_out0;
assign v_RD_5964_out0 = v_RD_7236_out0;
assign v_RD_5969_out0 = v_RD_7238_out0;
assign v_RD_5979_out0 = v_RD_7243_out0;
assign v_RD_6016_out0 = v_RD_7261_out0;
assign v_RD_6018_out0 = v_RD_7262_out0;
assign v_RD_6020_out0 = v_RD_7263_out0;
assign v_RD_6026_out0 = v_RD_7266_out0;
assign v_RD_6031_out0 = v_RD_7268_out0;
assign v_RD_6041_out0 = v_RD_7273_out0;
assign v_RD_6047_out0 = v_RD_7276_out0;
assign v_RD_6049_out0 = v_RD_7277_out0;
assign v_RD_6051_out0 = v_RD_7278_out0;
assign v_RD_6057_out0 = v_RD_7281_out0;
assign v_RD_6062_out0 = v_RD_7283_out0;
assign v_RD_6072_out0 = v_RD_7288_out0;
assign v_RD_6078_out0 = v_RD_7291_out0;
assign v_RD_6080_out0 = v_RD_7292_out0;
assign v_RD_6082_out0 = v_RD_7293_out0;
assign v_RD_6088_out0 = v_RD_7296_out0;
assign v_RD_6093_out0 = v_RD_7298_out0;
assign v_RD_6103_out0 = v_RD_7303_out0;
assign v_RD_6109_out0 = v_RD_7306_out0;
assign v_RD_6111_out0 = v_RD_7307_out0;
assign v_RD_6113_out0 = v_RD_7308_out0;
assign v_RD_6119_out0 = v_RD_7311_out0;
assign v_RD_6124_out0 = v_RD_7313_out0;
assign v_RD_6134_out0 = v_RD_7318_out0;
assign v_RD_6140_out0 = v_RD_7321_out0;
assign v_RD_6142_out0 = v_RD_7322_out0;
assign v_RD_6144_out0 = v_RD_7323_out0;
assign v_RD_6150_out0 = v_RD_7326_out0;
assign v_RD_6155_out0 = v_RD_7328_out0;
assign v_RD_6165_out0 = v_RD_7333_out0;
assign v_RD_6171_out0 = v_RD_7336_out0;
assign v_RD_6173_out0 = v_RD_7337_out0;
assign v_RD_6175_out0 = v_RD_7338_out0;
assign v_RD_6181_out0 = v_RD_7341_out0;
assign v_RD_6186_out0 = v_RD_7343_out0;
assign v_RD_6196_out0 = v_RD_7348_out0;
assign v_RD_6202_out0 = v_RD_7351_out0;
assign v_RD_6204_out0 = v_RD_7352_out0;
assign v_RD_6206_out0 = v_RD_7353_out0;
assign v_RD_6212_out0 = v_RD_7356_out0;
assign v_RD_6217_out0 = v_RD_7358_out0;
assign v_RD_6227_out0 = v_RD_7363_out0;
assign v_RD_6233_out0 = v_RD_7366_out0;
assign v_RD_6235_out0 = v_RD_7367_out0;
assign v_RD_6237_out0 = v_RD_7368_out0;
assign v_RD_6243_out0 = v_RD_7371_out0;
assign v_RD_6248_out0 = v_RD_7373_out0;
assign v_RD_6258_out0 = v_RD_7378_out0;
assign v_RD_6264_out0 = v_RD_7381_out0;
assign v_RD_6266_out0 = v_RD_7382_out0;
assign v_RD_6268_out0 = v_RD_7383_out0;
assign v_RD_6274_out0 = v_RD_7386_out0;
assign v_RD_6279_out0 = v_RD_7388_out0;
assign v_RD_6289_out0 = v_RD_7393_out0;
assign v_RD_6295_out0 = v_RD_7396_out0;
assign v_RD_6297_out0 = v_RD_7397_out0;
assign v_RD_6299_out0 = v_RD_7398_out0;
assign v_RD_6305_out0 = v_RD_7401_out0;
assign v_RD_6310_out0 = v_RD_7403_out0;
assign v_RD_6320_out0 = v_RD_7408_out0;
assign v_RD_6326_out0 = v_RD_7411_out0;
assign v_RD_6328_out0 = v_RD_7412_out0;
assign v_RD_6330_out0 = v_RD_7413_out0;
assign v_RD_6336_out0 = v_RD_7416_out0;
assign v_RD_6341_out0 = v_RD_7418_out0;
assign v_RD_6351_out0 = v_RD_7423_out0;
assign v_RD_6418_out0 = v_RD_7455_out0;
assign v_RD_6420_out0 = v_RD_7456_out0;
assign v_RD_6422_out0 = v_RD_7457_out0;
assign v_RD_6428_out0 = v_RD_7460_out0;
assign v_RD_6433_out0 = v_RD_7462_out0;
assign v_RD_6443_out0 = v_RD_7467_out0;
assign v_RD_6480_out0 = v_RD_7485_out0;
assign v_RD_6482_out0 = v_RD_7486_out0;
assign v_RD_6484_out0 = v_RD_7487_out0;
assign v_RD_6490_out0 = v_RD_7490_out0;
assign v_RD_6495_out0 = v_RD_7492_out0;
assign v_RD_6505_out0 = v_RD_7497_out0;
assign v_RD_6511_out0 = v_RD_7500_out0;
assign v_RD_6513_out0 = v_RD_7501_out0;
assign v_RD_6515_out0 = v_RD_7502_out0;
assign v_RD_6521_out0 = v_RD_7505_out0;
assign v_RD_6526_out0 = v_RD_7507_out0;
assign v_RD_6536_out0 = v_RD_7512_out0;
assign v_RD_6542_out0 = v_RD_7515_out0;
assign v_RD_6544_out0 = v_RD_7516_out0;
assign v_RD_6546_out0 = v_RD_7517_out0;
assign v_RD_6552_out0 = v_RD_7520_out0;
assign v_RD_6557_out0 = v_RD_7522_out0;
assign v_RD_6567_out0 = v_RD_7527_out0;
assign v_RD_6573_out0 = v_RD_7530_out0;
assign v_RD_6575_out0 = v_RD_7531_out0;
assign v_RD_6577_out0 = v_RD_7532_out0;
assign v_RD_6583_out0 = v_RD_7535_out0;
assign v_RD_6588_out0 = v_RD_7537_out0;
assign v_RD_6598_out0 = v_RD_7542_out0;
assign v_RD_6604_out0 = v_RD_7545_out0;
assign v_RD_6606_out0 = v_RD_7546_out0;
assign v_RD_6608_out0 = v_RD_7547_out0;
assign v_RD_6614_out0 = v_RD_7550_out0;
assign v_RD_6619_out0 = v_RD_7552_out0;
assign v_RD_6629_out0 = v_RD_7557_out0;
assign v_RD_6635_out0 = v_RD_7560_out0;
assign v_RD_6637_out0 = v_RD_7561_out0;
assign v_RD_6639_out0 = v_RD_7562_out0;
assign v_RD_6645_out0 = v_RD_7565_out0;
assign v_RD_6650_out0 = v_RD_7567_out0;
assign v_RD_6660_out0 = v_RD_7572_out0;
assign v_RD_6666_out0 = v_RD_7575_out0;
assign v_RD_6668_out0 = v_RD_7576_out0;
assign v_RD_6670_out0 = v_RD_7577_out0;
assign v_RD_6676_out0 = v_RD_7580_out0;
assign v_RD_6681_out0 = v_RD_7582_out0;
assign v_RD_6691_out0 = v_RD_7587_out0;
assign v_RD_6697_out0 = v_RD_7590_out0;
assign v_RD_6699_out0 = v_RD_7591_out0;
assign v_RD_6701_out0 = v_RD_7592_out0;
assign v_RD_6707_out0 = v_RD_7595_out0;
assign v_RD_6712_out0 = v_RD_7597_out0;
assign v_RD_6722_out0 = v_RD_7602_out0;
assign v_RD_6728_out0 = v_RD_7605_out0;
assign v_RD_6730_out0 = v_RD_7606_out0;
assign v_RD_6732_out0 = v_RD_7607_out0;
assign v_RD_6738_out0 = v_RD_7610_out0;
assign v_RD_6743_out0 = v_RD_7612_out0;
assign v_RD_6753_out0 = v_RD_7617_out0;
assign v_RD_6759_out0 = v_RD_7620_out0;
assign v_RD_6761_out0 = v_RD_7621_out0;
assign v_RD_6763_out0 = v_RD_7622_out0;
assign v_RD_6769_out0 = v_RD_7625_out0;
assign v_RD_6774_out0 = v_RD_7627_out0;
assign v_RD_6784_out0 = v_RD_7632_out0;
assign v_ADDER_IN_10995_out0 = v__10783_out0;
assign v_NOTUSED_325_out0 = v__3907_out0;
assign v_NOTUSED_326_out0 = v__3908_out0;
assign v_ANDOUT_630_out0 = v__1867_out0;
assign v_ANDOUT_632_out0 = v__1869_out0;
assign v__4483_out0 = v_MUX1_6_out0[1:0];
assign v__4483_out1 = v_MUX1_6_out0[15:14];
assign v__4484_out0 = v_MUX1_7_out0[1:0];
assign v__4484_out1 = v_MUX1_7_out0[15:14];
assign v__4591_out0 = { v__3907_out1,v_C1_8815_out0 };
assign v__4592_out0 = { v__3908_out1,v_C1_8816_out0 };
assign v__5846_out0 = v_A1_3174_out0[11:0];
assign v__5846_out1 = v_A1_3174_out0[15:4];
assign v__5847_out0 = v_A1_3175_out0[11:0];
assign v__5847_out1 = v_A1_3175_out0[15:4];
assign v_COUT_10547_out0 = v_A1_3174_out1;
assign v_COUT_10548_out0 = v_A1_3175_out1;
assign v_RMN_13437_out0 = v_A1_3174_out0;
assign v_RMN_13438_out0 = v_A1_3175_out0;
assign v_OUT1_1972_out0 = v__4591_out0;
assign v_OUT1_1973_out0 = v__4592_out0;
assign v_NOTUSE_2399_out0 = v__5846_out1;
assign v_NOTUSE_2400_out0 = v__5847_out1;
assign v__10910_out0 = v_ANDOUT_630_out0[0:0];
assign v__10910_out1 = v_ANDOUT_630_out0[15:15];
assign v__10911_out0 = v_ANDOUT_632_out0[0:0];
assign v__10911_out1 = v_ANDOUT_632_out0[15:15];
assign v_UNUSED_11244_out0 = v__4483_out0;
assign v_UNUSED_11245_out0 = v__4484_out0;
assign v__13482_out0 = { v__4483_out1,v_C1_6793_out0 };
assign v__13483_out0 = { v__4484_out1,v_C1_6794_out0 };
assign v_MUX2_13656_out0 = v_G6_13258_out0 ? v__5846_out0 : v__3035_out0;
assign v_MUX2_13657_out0 = v_G6_13259_out0 ? v__5847_out0 : v__3036_out0;
assign v_CIN_2356_out0 = v__10910_out1;
assign v_CIN_2371_out0 = v__10911_out1;
assign v_MUX2_10841_out0 = v_LSR_13331_out0 ? v__13482_out0 : v_MUX1_6_out0;
assign v_MUX2_10842_out0 = v_LSR_13332_out0 ? v__13483_out0 : v_MUX1_7_out0;
assign v_EA_13516_out0 = v_MUX2_13656_out0;
assign v_EA_13517_out0 = v_MUX2_13657_out0;
assign v_MUX5_13670_out0 = v_0_3022_out0 ? v_OUT1_1972_out0 : v_IN_13668_out0;
assign v_MUX5_13671_out0 = v_0_3023_out0 ? v_OUT1_1973_out0 : v_IN_13669_out0;
assign v__469_out0 = v_CIN_2356_out0[8:8];
assign v__484_out0 = v_CIN_2371_out0[8:8];
assign v__1774_out0 = v_CIN_2356_out0[6:6];
assign v__1789_out0 = v_CIN_2371_out0[6:6];
assign v_IN_1964_out0 = v_MUX2_10841_out0;
assign v_IN_1965_out0 = v_MUX2_10842_out0;
assign v__2156_out0 = v_CIN_2356_out0[3:3];
assign v__2171_out0 = v_CIN_2371_out0[3:3];
assign v_RAMADDRMUX_2232_out0 = v_EA_13516_out0;
assign v_RAMADDRMUX_2233_out0 = v_EA_13517_out0;
assign v__2503_out0 = v_CIN_2356_out0[0:0];
assign v__2518_out0 = v_CIN_2371_out0[0:0];
assign v__3052_out0 = v_CIN_2356_out0[9:9];
assign v__3067_out0 = v_CIN_2371_out0[9:9];
assign v__3086_out0 = v_CIN_2356_out0[2:2];
assign v__3101_out0 = v_CIN_2371_out0[2:2];
assign v__3140_out0 = v_CIN_2356_out0[7:7];
assign v__3155_out0 = v_CIN_2371_out0[7:7];
assign v__3824_out0 = v_CIN_2356_out0[1:1];
assign v__3839_out0 = v_CIN_2371_out0[1:1];
assign v__3862_out0 = v_CIN_2356_out0[10:10];
assign v__3877_out0 = v_CIN_2371_out0[10:10];
assign v__6801_out0 = v_CIN_2356_out0[11:11];
assign v__6816_out0 = v_CIN_2371_out0[11:11];
assign v__7645_out0 = v_CIN_2356_out0[12:12];
assign v__7660_out0 = v_CIN_2371_out0[12:12];
assign v__8700_out0 = v_CIN_2356_out0[13:13];
assign v__8715_out0 = v_CIN_2371_out0[13:13];
assign v__8770_out0 = v_CIN_2356_out0[14:14];
assign v__8785_out0 = v_CIN_2371_out0[14:14];
assign v__10720_out0 = v_CIN_2356_out0[5:5];
assign v__10735_out0 = v_CIN_2371_out0[5:5];
assign v_IN1_10992_out0 = v_MUX5_13670_out0;
assign v_IN1_10993_out0 = v_MUX5_13671_out0;
assign v__13449_out0 = v_CIN_2356_out0[4:4];
assign v__13464_out0 = v_CIN_2371_out0[4:4];
assign v_RAMADDRMUX_92_out0 = v_RAMADDRMUX_2232_out0;
assign v_RAMADDRMUX_93_out0 = v_RAMADDRMUX_2233_out0;
assign v__627_out0 = v_IN_1964_out0[1:0];
assign v__627_out1 = v_IN_1964_out0[15:14];
assign v__628_out0 = v_IN_1965_out0[1:0];
assign v__628_out1 = v_IN_1965_out0[15:14];
assign v_RM_3370_out0 = v__7645_out0;
assign v_RM_3371_out0 = v__8770_out0;
assign v_RM_3372_out0 = v__10720_out0;
assign v_RM_3373_out0 = v__13449_out0;
assign v_RM_3374_out0 = v__8700_out0;
assign v_RM_3375_out0 = v__3052_out0;
assign v_RM_3376_out0 = v__3862_out0;
assign v_RM_3377_out0 = v__3824_out0;
assign v_RM_3378_out0 = v__2156_out0;
assign v_RM_3379_out0 = v__1774_out0;
assign v_RM_3380_out0 = v__3140_out0;
assign v_RM_3381_out0 = v__6801_out0;
assign v_RM_3382_out0 = v__469_out0;
assign v_RM_3383_out0 = v__3086_out0;
assign v_RM_3594_out0 = v__7660_out0;
assign v_RM_3595_out0 = v__8785_out0;
assign v_RM_3596_out0 = v__10735_out0;
assign v_RM_3597_out0 = v__13464_out0;
assign v_RM_3598_out0 = v__8715_out0;
assign v_RM_3599_out0 = v__3067_out0;
assign v_RM_3600_out0 = v__3877_out0;
assign v_RM_3601_out0 = v__3839_out0;
assign v_RM_3602_out0 = v__2171_out0;
assign v_RM_3603_out0 = v__1789_out0;
assign v_RM_3604_out0 = v__3155_out0;
assign v_RM_3605_out0 = v__6816_out0;
assign v_RM_3606_out0 = v__484_out0;
assign v_RM_3607_out0 = v__3101_out0;
assign v__10823_out0 = v_IN_1964_out0[15:15];
assign v__10824_out0 = v_IN_1965_out0[15:15];
assign v_RM_11343_out0 = v__2503_out0;
assign v_RM_11807_out0 = v__2518_out0;
assign v__13550_out0 = v_IN1_10992_out0[1:0];
assign v__13550_out1 = v_IN1_10992_out0[10:9];
assign v__13551_out0 = v_IN1_10993_out0[1:0];
assign v__13551_out1 = v_IN1_10993_out0[10:9];
assign v_NOTUSED_445_out0 = v__13550_out0;
assign v_NOTUSED_446_out0 = v__13551_out0;
assign v_NOTUSED_447_out0 = v__627_out0;
assign v_NOTUSED_448_out0 = v__628_out0;
assign v_G1_7758_out0 = ((v_RD_5903_out0 && !v_RM_11343_out0) || (!v_RD_5903_out0) && v_RM_11343_out0);
assign v_G1_8222_out0 = ((v_RD_6367_out0 && !v_RM_11807_out0) || (!v_RD_6367_out0) && v_RM_11807_out0);
assign v__10354_out0 = { v__627_out1,v__10823_out0 };
assign v__10355_out0 = { v__628_out1,v__10824_out0 };
assign v_RAMADDRMUX_10542_out0 = v_RAMADDRMUX_92_out0;
assign v_RAMADDRMUX_10543_out0 = v_RAMADDRMUX_93_out0;
assign v_RM_11333_out0 = v_RM_3370_out0;
assign v_RM_11335_out0 = v_RM_3371_out0;
assign v_RM_11337_out0 = v_RM_3372_out0;
assign v_RM_11339_out0 = v_RM_3373_out0;
assign v_RM_11341_out0 = v_RM_3374_out0;
assign v_RM_11345_out0 = v_RM_3375_out0;
assign v_RM_11347_out0 = v_RM_3376_out0;
assign v_RM_11349_out0 = v_RM_3377_out0;
assign v_RM_11351_out0 = v_RM_3378_out0;
assign v_RM_11353_out0 = v_RM_3379_out0;
assign v_RM_11355_out0 = v_RM_3380_out0;
assign v_RM_11357_out0 = v_RM_3381_out0;
assign v_RM_11359_out0 = v_RM_3382_out0;
assign v_RM_11361_out0 = v_RM_3383_out0;
assign v_RM_11797_out0 = v_RM_3594_out0;
assign v_RM_11799_out0 = v_RM_3595_out0;
assign v_RM_11801_out0 = v_RM_3596_out0;
assign v_RM_11803_out0 = v_RM_3597_out0;
assign v_RM_11805_out0 = v_RM_3598_out0;
assign v_RM_11809_out0 = v_RM_3599_out0;
assign v_RM_11811_out0 = v_RM_3600_out0;
assign v_RM_11813_out0 = v_RM_3601_out0;
assign v_RM_11815_out0 = v_RM_3602_out0;
assign v_RM_11817_out0 = v_RM_3603_out0;
assign v_RM_11819_out0 = v_RM_3604_out0;
assign v_RM_11821_out0 = v_RM_3605_out0;
assign v_RM_11823_out0 = v_RM_3606_out0;
assign v_RM_11825_out0 = v_RM_3607_out0;
assign v_G2_12294_out0 = v_RD_5903_out0 && v_RM_11343_out0;
assign v_G2_12758_out0 = v_RD_6367_out0 && v_RM_11807_out0;
assign v__13761_out0 = { v__13550_out1,v_C1_3205_out0 };
assign v__13762_out0 = { v__13551_out1,v_C1_3206_out0 };
assign v__1172_out0 = { v__10354_out0,v__10823_out0 };
assign v__1173_out0 = { v__10355_out0,v__10824_out0 };
assign v_OUT1_3853_out0 = v__13761_out0;
assign v_OUT1_3854_out0 = v__13762_out0;
assign v_CARRY_4903_out0 = v_G2_12294_out0;
assign v_CARRY_5367_out0 = v_G2_12758_out0;
assign v_G1_7748_out0 = ((v_RD_5893_out0 && !v_RM_11333_out0) || (!v_RD_5893_out0) && v_RM_11333_out0);
assign v_G1_7750_out0 = ((v_RD_5895_out0 && !v_RM_11335_out0) || (!v_RD_5895_out0) && v_RM_11335_out0);
assign v_G1_7752_out0 = ((v_RD_5897_out0 && !v_RM_11337_out0) || (!v_RD_5897_out0) && v_RM_11337_out0);
assign v_G1_7754_out0 = ((v_RD_5899_out0 && !v_RM_11339_out0) || (!v_RD_5899_out0) && v_RM_11339_out0);
assign v_G1_7756_out0 = ((v_RD_5901_out0 && !v_RM_11341_out0) || (!v_RD_5901_out0) && v_RM_11341_out0);
assign v_G1_7760_out0 = ((v_RD_5905_out0 && !v_RM_11345_out0) || (!v_RD_5905_out0) && v_RM_11345_out0);
assign v_G1_7762_out0 = ((v_RD_5907_out0 && !v_RM_11347_out0) || (!v_RD_5907_out0) && v_RM_11347_out0);
assign v_G1_7764_out0 = ((v_RD_5909_out0 && !v_RM_11349_out0) || (!v_RD_5909_out0) && v_RM_11349_out0);
assign v_G1_7766_out0 = ((v_RD_5911_out0 && !v_RM_11351_out0) || (!v_RD_5911_out0) && v_RM_11351_out0);
assign v_G1_7768_out0 = ((v_RD_5913_out0 && !v_RM_11353_out0) || (!v_RD_5913_out0) && v_RM_11353_out0);
assign v_G1_7770_out0 = ((v_RD_5915_out0 && !v_RM_11355_out0) || (!v_RD_5915_out0) && v_RM_11355_out0);
assign v_G1_7772_out0 = ((v_RD_5917_out0 && !v_RM_11357_out0) || (!v_RD_5917_out0) && v_RM_11357_out0);
assign v_G1_7774_out0 = ((v_RD_5919_out0 && !v_RM_11359_out0) || (!v_RD_5919_out0) && v_RM_11359_out0);
assign v_G1_7776_out0 = ((v_RD_5921_out0 && !v_RM_11361_out0) || (!v_RD_5921_out0) && v_RM_11361_out0);
assign v_G1_8212_out0 = ((v_RD_6357_out0 && !v_RM_11797_out0) || (!v_RD_6357_out0) && v_RM_11797_out0);
assign v_G1_8214_out0 = ((v_RD_6359_out0 && !v_RM_11799_out0) || (!v_RD_6359_out0) && v_RM_11799_out0);
assign v_G1_8216_out0 = ((v_RD_6361_out0 && !v_RM_11801_out0) || (!v_RD_6361_out0) && v_RM_11801_out0);
assign v_G1_8218_out0 = ((v_RD_6363_out0 && !v_RM_11803_out0) || (!v_RD_6363_out0) && v_RM_11803_out0);
assign v_G1_8220_out0 = ((v_RD_6365_out0 && !v_RM_11805_out0) || (!v_RD_6365_out0) && v_RM_11805_out0);
assign v_G1_8224_out0 = ((v_RD_6369_out0 && !v_RM_11809_out0) || (!v_RD_6369_out0) && v_RM_11809_out0);
assign v_G1_8226_out0 = ((v_RD_6371_out0 && !v_RM_11811_out0) || (!v_RD_6371_out0) && v_RM_11811_out0);
assign v_G1_8228_out0 = ((v_RD_6373_out0 && !v_RM_11813_out0) || (!v_RD_6373_out0) && v_RM_11813_out0);
assign v_G1_8230_out0 = ((v_RD_6375_out0 && !v_RM_11815_out0) || (!v_RD_6375_out0) && v_RM_11815_out0);
assign v_G1_8232_out0 = ((v_RD_6377_out0 && !v_RM_11817_out0) || (!v_RD_6377_out0) && v_RM_11817_out0);
assign v_G1_8234_out0 = ((v_RD_6379_out0 && !v_RM_11819_out0) || (!v_RD_6379_out0) && v_RM_11819_out0);
assign v_G1_8236_out0 = ((v_RD_6381_out0 && !v_RM_11821_out0) || (!v_RD_6381_out0) && v_RM_11821_out0);
assign v_G1_8238_out0 = ((v_RD_6383_out0 && !v_RM_11823_out0) || (!v_RD_6383_out0) && v_RM_11823_out0);
assign v_G1_8240_out0 = ((v_RD_6385_out0 && !v_RM_11825_out0) || (!v_RD_6385_out0) && v_RM_11825_out0);
assign v_RAM_ADDRESS_MUX_8803_out0 = v_RAMADDRMUX_10542_out0;
assign v_RAM_ADDRESS_MUX_8804_out0 = v_RAMADDRMUX_10543_out0;
assign v_S_8904_out0 = v_G1_7758_out0;
assign v_S_9368_out0 = v_G1_8222_out0;
assign v_G2_12284_out0 = v_RD_5893_out0 && v_RM_11333_out0;
assign v_G2_12286_out0 = v_RD_5895_out0 && v_RM_11335_out0;
assign v_G2_12288_out0 = v_RD_5897_out0 && v_RM_11337_out0;
assign v_G2_12290_out0 = v_RD_5899_out0 && v_RM_11339_out0;
assign v_G2_12292_out0 = v_RD_5901_out0 && v_RM_11341_out0;
assign v_G2_12296_out0 = v_RD_5905_out0 && v_RM_11345_out0;
assign v_G2_12298_out0 = v_RD_5907_out0 && v_RM_11347_out0;
assign v_G2_12300_out0 = v_RD_5909_out0 && v_RM_11349_out0;
assign v_G2_12302_out0 = v_RD_5911_out0 && v_RM_11351_out0;
assign v_G2_12304_out0 = v_RD_5913_out0 && v_RM_11353_out0;
assign v_G2_12306_out0 = v_RD_5915_out0 && v_RM_11355_out0;
assign v_G2_12308_out0 = v_RD_5917_out0 && v_RM_11357_out0;
assign v_G2_12310_out0 = v_RD_5919_out0 && v_RM_11359_out0;
assign v_G2_12312_out0 = v_RD_5921_out0 && v_RM_11361_out0;
assign v_G2_12748_out0 = v_RD_6357_out0 && v_RM_11797_out0;
assign v_G2_12750_out0 = v_RD_6359_out0 && v_RM_11799_out0;
assign v_G2_12752_out0 = v_RD_6361_out0 && v_RM_11801_out0;
assign v_G2_12754_out0 = v_RD_6363_out0 && v_RM_11803_out0;
assign v_G2_12756_out0 = v_RD_6365_out0 && v_RM_11805_out0;
assign v_G2_12760_out0 = v_RD_6369_out0 && v_RM_11809_out0;
assign v_G2_12762_out0 = v_RD_6371_out0 && v_RM_11811_out0;
assign v_G2_12764_out0 = v_RD_6373_out0 && v_RM_11813_out0;
assign v_G2_12766_out0 = v_RD_6375_out0 && v_RM_11815_out0;
assign v_G2_12768_out0 = v_RD_6377_out0 && v_RM_11817_out0;
assign v_G2_12770_out0 = v_RD_6379_out0 && v_RM_11819_out0;
assign v_G2_12772_out0 = v_RD_6381_out0 && v_RM_11821_out0;
assign v_G2_12774_out0 = v_RD_6383_out0 && v_RM_11823_out0;
assign v_G2_12776_out0 = v_RD_6385_out0 && v_RM_11825_out0;
assign v_RAM_ADDRES_MUX_13649_out0 = v_RAMADDRMUX_10542_out0;
assign v_RAM_ADDRES_MUX_13650_out0 = v_RAMADDRMUX_10543_out0;
assign v_MUX4_552_out0 = v_1_3817_out0 ? v_OUT1_3853_out0 : v_MUX5_13670_out0;
assign v_MUX4_553_out0 = v_1_3818_out0 ? v_OUT1_3854_out0 : v_MUX5_13671_out0;
assign v_ADRESS1_1906_out0 = v_RAM_ADDRES_MUX_13649_out0;
assign v_S_4666_out0 = v_S_8904_out0;
assign v_S_4681_out0 = v_S_9368_out0;
assign v_CARRY_4893_out0 = v_G2_12284_out0;
assign v_CARRY_4895_out0 = v_G2_12286_out0;
assign v_CARRY_4897_out0 = v_G2_12288_out0;
assign v_CARRY_4899_out0 = v_G2_12290_out0;
assign v_CARRY_4901_out0 = v_G2_12292_out0;
assign v_CARRY_4905_out0 = v_G2_12296_out0;
assign v_CARRY_4907_out0 = v_G2_12298_out0;
assign v_CARRY_4909_out0 = v_G2_12300_out0;
assign v_CARRY_4911_out0 = v_G2_12302_out0;
assign v_CARRY_4913_out0 = v_G2_12304_out0;
assign v_CARRY_4915_out0 = v_G2_12306_out0;
assign v_CARRY_4917_out0 = v_G2_12308_out0;
assign v_CARRY_4919_out0 = v_G2_12310_out0;
assign v_CARRY_4921_out0 = v_G2_12312_out0;
assign v_CARRY_5357_out0 = v_G2_12748_out0;
assign v_CARRY_5359_out0 = v_G2_12750_out0;
assign v_CARRY_5361_out0 = v_G2_12752_out0;
assign v_CARRY_5363_out0 = v_G2_12754_out0;
assign v_CARRY_5365_out0 = v_G2_12756_out0;
assign v_CARRY_5369_out0 = v_G2_12760_out0;
assign v_CARRY_5371_out0 = v_G2_12762_out0;
assign v_CARRY_5373_out0 = v_G2_12764_out0;
assign v_CARRY_5375_out0 = v_G2_12766_out0;
assign v_CARRY_5377_out0 = v_G2_12768_out0;
assign v_CARRY_5379_out0 = v_G2_12770_out0;
assign v_CARRY_5381_out0 = v_G2_12772_out0;
assign v_CARRY_5383_out0 = v_G2_12774_out0;
assign v_CARRY_5385_out0 = v_G2_12776_out0;
assign v_RAMADDRMUX_7066_out0 = v_RAM_ADDRESS_MUX_8803_out0;
assign v_RAMADDRMUX_7067_out0 = v_RAM_ADDRESS_MUX_8804_out0;
assign v_OUT_8852_out0 = v__1172_out0;
assign v_OUT_8853_out0 = v__1173_out0;
assign v_S_8894_out0 = v_G1_7748_out0;
assign v_S_8896_out0 = v_G1_7750_out0;
assign v_S_8898_out0 = v_G1_7752_out0;
assign v_S_8900_out0 = v_G1_7754_out0;
assign v_S_8902_out0 = v_G1_7756_out0;
assign v_S_8906_out0 = v_G1_7760_out0;
assign v_S_8908_out0 = v_G1_7762_out0;
assign v_S_8910_out0 = v_G1_7764_out0;
assign v_S_8912_out0 = v_G1_7766_out0;
assign v_S_8914_out0 = v_G1_7768_out0;
assign v_S_8916_out0 = v_G1_7770_out0;
assign v_S_8918_out0 = v_G1_7772_out0;
assign v_S_8920_out0 = v_G1_7774_out0;
assign v_S_8922_out0 = v_G1_7776_out0;
assign v_S_9358_out0 = v_G1_8212_out0;
assign v_S_9360_out0 = v_G1_8214_out0;
assign v_S_9362_out0 = v_G1_8216_out0;
assign v_S_9364_out0 = v_G1_8218_out0;
assign v_S_9366_out0 = v_G1_8220_out0;
assign v_S_9370_out0 = v_G1_8224_out0;
assign v_S_9372_out0 = v_G1_8226_out0;
assign v_S_9374_out0 = v_G1_8228_out0;
assign v_S_9376_out0 = v_G1_8230_out0;
assign v_S_9378_out0 = v_G1_8232_out0;
assign v_S_9380_out0 = v_G1_8234_out0;
assign v_S_9382_out0 = v_G1_8236_out0;
assign v_S_9384_out0 = v_G1_8238_out0;
assign v_S_9386_out0 = v_G1_8240_out0;
assign v_CIN_9830_out0 = v_CARRY_4903_out0;
assign v_CIN_10054_out0 = v_CARRY_5367_out0;
assign v_ADRESS0_11217_out0 = v_RAM_ADDRES_MUX_13650_out0;
assign v__2437_out0 = v_RAMADDRMUX_7066_out0[3:0];
assign v__2437_out1 = v_RAMADDRMUX_7066_out0[11:8];
assign v__2438_out0 = v_RAMADDRMUX_7067_out0[3:0];
assign v__2438_out1 = v_RAMADDRMUX_7067_out0[11:8];
assign v_IN1_2848_out0 = v_MUX4_552_out0;
assign v_IN1_2849_out0 = v_MUX4_553_out0;
assign v_ADDRESS1_2854_out0 = v_ADRESS1_1906_out0;
assign v_MUX3_3133_out0 = v_ASR_13713_out0 ? v_OUT_8852_out0 : v_MUX2_10841_out0;
assign v_MUX3_3134_out0 = v_ASR_13714_out0 ? v_OUT_8853_out0 : v_MUX2_10842_out0;
assign v__3223_out0 = { v__10910_out0,v_S_4666_out0 };
assign v__3224_out0 = { v__10911_out0,v_S_4681_out0 };
assign v_EQ11_4465_out0 = v_RAMADDRMUX_7066_out0 == 12'h800;
assign v_EQ11_4466_out0 = v_RAMADDRMUX_7067_out0 == 12'h800;
assign v_RD_5910_out0 = v_CIN_9830_out0;
assign v_RD_6374_out0 = v_CIN_10054_out0;
assign v_ADDRESS0_10982_out0 = v_ADRESS0_11217_out0;
assign v_RM_11334_out0 = v_S_8894_out0;
assign v_RM_11336_out0 = v_S_8896_out0;
assign v_RM_11338_out0 = v_S_8898_out0;
assign v_RM_11340_out0 = v_S_8900_out0;
assign v_RM_11342_out0 = v_S_8902_out0;
assign v_RM_11346_out0 = v_S_8906_out0;
assign v_RM_11348_out0 = v_S_8908_out0;
assign v_RM_11350_out0 = v_S_8910_out0;
assign v_RM_11352_out0 = v_S_8912_out0;
assign v_RM_11354_out0 = v_S_8914_out0;
assign v_RM_11356_out0 = v_S_8916_out0;
assign v_RM_11358_out0 = v_S_8918_out0;
assign v_RM_11360_out0 = v_S_8920_out0;
assign v_RM_11362_out0 = v_S_8922_out0;
assign v_RM_11798_out0 = v_S_9358_out0;
assign v_RM_11800_out0 = v_S_9360_out0;
assign v_RM_11802_out0 = v_S_9362_out0;
assign v_RM_11804_out0 = v_S_9364_out0;
assign v_RM_11806_out0 = v_S_9366_out0;
assign v_RM_11810_out0 = v_S_9370_out0;
assign v_RM_11812_out0 = v_S_9372_out0;
assign v_RM_11814_out0 = v_S_9374_out0;
assign v_RM_11816_out0 = v_S_9376_out0;
assign v_RM_11818_out0 = v_S_9378_out0;
assign v_RM_11820_out0 = v_S_9380_out0;
assign v_RM_11822_out0 = v_S_9382_out0;
assign v_RM_11824_out0 = v_S_9384_out0;
assign v_RM_11826_out0 = v_S_9386_out0;
assign v__4703_out0 = v_IN1_2848_out0[3:0];
assign v__4703_out1 = v_IN1_2848_out0[10:7];
assign v__4704_out0 = v_IN1_2849_out0[3:0];
assign v__4704_out1 = v_IN1_2849_out0[10:7];
assign v__4816_out0 = v_MUX3_3133_out0[1:0];
assign v__4816_out1 = v_MUX3_3133_out0[15:14];
assign v__4817_out0 = v_MUX3_3134_out0[1:0];
assign v__4817_out1 = v_MUX3_3134_out0[15:14];
assign v_MUX1_7097_out0 = v_MUX_ENABLE_2349_out0 ? v_ADDRESS0_10982_out0 : v_ADDRESS1_2854_out0;
assign v_G1_7765_out0 = ((v_RD_5910_out0 && !v_RM_11350_out0) || (!v_RD_5910_out0) && v_RM_11350_out0);
assign v_G1_8229_out0 = ((v_RD_6374_out0 && !v_RM_11814_out0) || (!v_RD_6374_out0) && v_RM_11814_out0);
assign v_G2_12301_out0 = v_RD_5910_out0 && v_RM_11350_out0;
assign v_G2_12765_out0 = v_RD_6374_out0 && v_RM_11814_out0;
assign v__13317_out0 = v__2437_out1[3:0];
assign v__13317_out1 = v__2437_out1[7:4];
assign v__13318_out0 = v__2438_out1[3:0];
assign v__13318_out1 = v__2438_out1[7:4];
assign v_RAM_ADD_BYTE0_13382_out0 = v__2437_out0;
assign v_RAM_ADD_BYTE0_13383_out0 = v__2438_out0;
assign v_G22_13707_out0 = v_EQ11_4465_out0 && v_UART_11128_out0;
assign v_G22_13708_out0 = v_EQ11_4466_out0 && v_UART_11129_out0;
assign v__1209_out0 = { v__4816_out1,v__4816_out0 };
assign v__1210_out0 = { v__4817_out1,v__4817_out0 };
assign v_EQ1_2675_out0 = v__13317_out0 == 4'h1;
assign v_EQ1_2676_out0 = v__13318_out0 == 4'h1;
assign v__2971_out0 = { v__4703_out1,v_C1_10305_out0 };
assign v__2972_out0 = { v__4704_out1,v_C1_10306_out0 };
assign v_ADDRESS_4662_out0 = v_MUX1_7097_out0;
assign v_EQ9_4842_out0 = v_RAM_ADD_BYTE0_13382_out0 == 4'h2;
assign v_EQ9_4843_out0 = v_RAM_ADD_BYTE0_13383_out0 == 4'h2;
assign v_CARRY_4910_out0 = v_G2_12301_out0;
assign v_CARRY_5374_out0 = v_G2_12765_out0;
assign v_S_8911_out0 = v_G1_7765_out0;
assign v_S_9375_out0 = v_G1_8229_out0;
assign v_G23_10439_out0 = v_G22_13707_out0 && v_LOAD_3949_out0;
assign v_G23_10440_out0 = v_G22_13708_out0 && v_LOAD_3950_out0;
assign v_EQ01_10510_out0 = v_RAM_ADD_BYTE0_13382_out0 == 4'h1;
assign v_EQ01_10511_out0 = v_RAM_ADD_BYTE0_13383_out0 == 4'h1;
assign v_NOTUSED_10540_out0 = v__4703_out0;
assign v_NOTUSED_10541_out0 = v__4704_out0;
assign v_EQ8_10804_out0 = v__13317_out1 == 4'h8;
assign v_EQ8_10805_out0 = v__13318_out1 == 4'h8;
assign v_S_1241_out0 = v_S_8911_out0;
assign v_S_1465_out0 = v_S_9375_out0;
assign v_OUT1_1873_out0 = v__2971_out0;
assign v_OUT1_1874_out0 = v__2972_out0;
assign v_BYTE1_comp1_2443_out0 = v_EQ1_2675_out0;
assign v_BYTE1_comp1_2444_out0 = v_EQ1_2676_out0;
assign v_STAT_INSTRUCTION_2855_out0 = v_G23_10439_out0;
assign v_STAT_INSTRUCTION_2856_out0 = v_G23_10440_out0;
assign v_G1_4017_out0 = v_CARRY_4910_out0 || v_CARRY_4909_out0;
assign v_G1_4241_out0 = v_CARRY_5374_out0 || v_CARRY_5373_out0;
assign v_BYTE2_COMP8_7695_out0 = v_EQ8_10804_out0;
assign v_BYTE2_COMP8_7696_out0 = v_EQ8_10805_out0;
assign v_ADRESS_8683_out0 = v_ADDRESS_4662_out0;
assign v_MUX4_10524_out0 = v_ROR_3286_out0 ? v__1209_out0 : v_MUX3_3133_out0;
assign v_MUX4_10525_out0 = v_ROR_3287_out0 ? v__1210_out0 : v_MUX3_3134_out0;
assign v_COUT_709_out0 = v_G1_4017_out0;
assign v_COUT_933_out0 = v_G1_4241_out0;
assign v_MUX5_1185_out0 = v_EN_10474_out0 ? v_MUX4_10524_out0 : v_IN_8838_out0;
assign v_MUX5_1186_out0 = v_EN_10475_out0 ? v_MUX4_10525_out0 : v_IN_8839_out0;
assign v_STAT_INSTRUCTION_2434_out0 = v_STAT_INSTRUCTION_2855_out0;
assign v_STAT_INSTRUCTION_2435_out0 = v_STAT_INSTRUCTION_2856_out0;
assign v_G2_3245_out0 = v_EQ01_10510_out0 && v_BYTE2_COMP8_7695_out0;
assign v_G2_3246_out0 = v_EQ01_10511_out0 && v_BYTE2_COMP8_7696_out0;
assign v_BYTE_COMP1_3262_out0 = v_BYTE1_comp1_2443_out0;
assign v_BYTE_COMP1_3263_out0 = v_BYTE1_comp1_2444_out0;
assign v_G20_11147_out0 = v_BYTE2_COMP8_7695_out0 && v_EQ9_4842_out0;
assign v_G20_11148_out0 = v_BYTE2_COMP8_7696_out0 && v_EQ9_4843_out0;
assign v_MUX3_13312_out0 = v_2_1763_out0 ? v_OUT1_1873_out0 : v_MUX4_552_out0;
assign v_MUX3_13313_out0 = v_2_1764_out0 ? v_OUT1_1874_out0 : v_MUX4_553_out0;
assign v_MUX3_13335_out0 = v_BYTE1_comp1_2443_out0 ? v__9791_out0 : v__7081_out0;
assign v_MUX3_13336_out0 = v_BYTE1_comp1_2444_out0 ? v__9792_out0 : v__7082_out0;
assign v_BYTE_COMP1_9796_out0 = v_BYTE_COMP1_3262_out0;
assign v_BYTE_COMP1_9797_out0 = v_BYTE_COMP1_3263_out0;
assign v_CIN_9836_out0 = v_COUT_709_out0;
assign v_CIN_10060_out0 = v_COUT_933_out0;
assign v_STAT_INSTRUCTION_10272_out0 = v_STAT_INSTRUCTION_2434_out0;
assign v_STAT_INSTRUCTION_10273_out0 = v_STAT_INSTRUCTION_2435_out0;
assign v_G14_10407_out0 = v_G2_3245_out0 && v_UART_11128_out0;
assign v_G14_10408_out0 = v_G2_3246_out0 && v_UART_11129_out0;
assign v_G18_11204_out0 = v_G20_11147_out0 && v_UART_11128_out0;
assign v_G18_11205_out0 = v_G20_11148_out0 && v_UART_11129_out0;
assign v_OUT_12236_out0 = v_MUX5_1185_out0;
assign v_OUT_12237_out0 = v_MUX5_1186_out0;
assign v_IN1_13711_out0 = v_MUX3_13312_out0;
assign v_IN1_13712_out0 = v_MUX3_13313_out0;
assign v_byte_comp_10_2318_out0 = v_BYTE_COMP1_9797_out0;
assign v_byte_comp_11_2645_out0 = v_BYTE_COMP1_9796_out0;
assign v_IN_2664_out0 = v_OUT_12236_out0;
assign v_IN_2665_out0 = v_OUT_12237_out0;
assign v__2680_out0 = v_IN1_13711_out0[7:0];
assign v__2680_out1 = v_IN1_13711_out0[10:3];
assign v__2681_out0 = v_IN1_13712_out0[7:0];
assign v__2681_out1 = v_IN1_13712_out0[10:3];
assign v_G19_4663_out0 = v_G18_11204_out0 && v_STORE_221_out0;
assign v_G19_4664_out0 = v_G18_11205_out0 && v_STORE_222_out0;
assign v_RD_5922_out0 = v_CIN_9836_out0;
assign v_RD_6386_out0 = v_CIN_10060_out0;
assign v_G16_13388_out0 = v_G14_10407_out0 && v_LOAD_3949_out0;
assign v_G16_13389_out0 = v_G14_10408_out0 && v_LOAD_3950_out0;
assign v_NOTUSED_683_out0 = v__2680_out0;
assign v_NOTUSED_684_out0 = v__2681_out0;
assign v_BYTE_COMP_11_1163_out0 = v_byte_comp_11_2645_out0;
assign v__2411_out0 = v_IN_2664_out0[11:0];
assign v__2411_out1 = v_IN_2664_out0[15:4];
assign v__2412_out0 = v_IN_2665_out0[11:0];
assign v__2412_out1 = v_IN_2665_out0[15:4];
assign v_G21_2885_out0 = v_G19_4663_out0 && v_EXEC1_3038_out0;
assign v_G21_2886_out0 = v_G19_4664_out0 && v_EXEC1_3039_out0;
assign v_G1_7777_out0 = ((v_RD_5922_out0 && !v_RM_11362_out0) || (!v_RD_5922_out0) && v_RM_11362_out0);
assign v_G1_8241_out0 = ((v_RD_6386_out0 && !v_RM_11826_out0) || (!v_RD_6386_out0) && v_RM_11826_out0);
assign v_RX_INSTRUCTION_11170_out0 = v_G16_13388_out0;
assign v_RX_INSTRUCTION_11171_out0 = v_G16_13389_out0;
assign v_G2_12313_out0 = v_RD_5922_out0 && v_RM_11362_out0;
assign v_G2_12777_out0 = v_RD_6386_out0 && v_RM_11826_out0;
assign v__13484_out0 = { v__2680_out1,v_C1_10266_out0 };
assign v__13485_out0 = { v__2681_out1,v_C1_10267_out0 };
assign v_IN_13548_out0 = v_IN_2664_out0;
assign v_IN_13549_out0 = v_IN_2665_out0;
assign v_BYTE_COMP_10_13611_out0 = v_byte_comp_10_2318_out0;
assign v_TX_INSTRUCTION_62_out0 = v_G21_2885_out0;
assign v_TX_INSTRUCTION_63_out0 = v_G21_2886_out0;
assign v_RX_INSTRUCTION_94_out0 = v_RX_INSTRUCTION_11170_out0;
assign v_RX_INSTRUCTION_95_out0 = v_RX_INSTRUCTION_11171_out0;
assign v_NOTUSED1_1897_out0 = v__2411_out1;
assign v_NOTUSED1_1898_out0 = v__2412_out1;
assign v__2678_out0 = { v_C1_6919_out0,v__2411_out0 };
assign v__2679_out0 = { v_C1_6920_out0,v__2412_out0 };
assign v_OUT1_3294_out0 = v__13484_out0;
assign v_OUT1_3295_out0 = v__13485_out0;
assign v_CARRY_4922_out0 = v_G2_12313_out0;
assign v_CARRY_5386_out0 = v_G2_12777_out0;
assign v_S_8923_out0 = v_G1_7777_out0;
assign v_S_9387_out0 = v_G1_8241_out0;
assign v_MUX1_11141_out0 = v_RX_INSTRUCTION_11170_out0 ? v_MUX3_13335_out0 : v_RAM_OUT_11214_out0;
assign v_MUX1_11142_out0 = v_RX_INSTRUCTION_11171_out0 ? v_MUX3_13336_out0 : v_RAM_OUT_11215_out0;
assign v_S_1247_out0 = v_S_8923_out0;
assign v_S_1471_out0 = v_S_9387_out0;
assign v_RX_INSTRUCTION_3258_out0 = v_RX_INSTRUCTION_94_out0;
assign v_RX_INSTRUCTION_3259_out0 = v_RX_INSTRUCTION_95_out0;
assign v_G1_4023_out0 = v_CARRY_4922_out0 || v_CARRY_4921_out0;
assign v_G1_4247_out0 = v_CARRY_5386_out0 || v_CARRY_5385_out0;
assign v_MUX1_4844_out0 = v_LSL_3047_out0 ? v__2678_out0 : v_IN_13548_out0;
assign v_MUX1_4845_out0 = v_LSL_3048_out0 ? v__2679_out0 : v_IN_13549_out0;
assign v_TX_INSTRUCTION_7012_out0 = v_TX_INSTRUCTION_62_out0;
assign v_TX_INSTRUCTION_7013_out0 = v_TX_INSTRUCTION_63_out0;
assign v_MUX1_7143_out0 = v_3_13619_out0 ? v_OUT1_3294_out0 : v_MUX3_13312_out0;
assign v_MUX1_7144_out0 = v_3_13620_out0 ? v_OUT1_3295_out0 : v_MUX3_13313_out0;
assign v_REGISTER_INPUT_13270_out0 = v_MUX1_11141_out0;
assign v_REGISTER_INPUT_13271_out0 = v_MUX1_11142_out0;
assign v_COUT_715_out0 = v_G1_4023_out0;
assign v_COUT_939_out0 = v_G1_4247_out0;
assign v_RX_INSTRUCTION_2343_out0 = v_RX_INSTRUCTION_3258_out0;
assign v_RX_INSTRUCTION_2344_out0 = v_RX_INSTRUCTION_3259_out0;
assign v_shifted1_2666_out0 = v_MUX1_7143_out0;
assign v_shifted1_2667_out0 = v_MUX1_7144_out0;
assign v_REGISTE_IN_4490_out0 = v_REGISTER_INPUT_13270_out0;
assign v_REGISTE_IN_4491_out0 = v_REGISTER_INPUT_13271_out0;
assign v__4585_out0 = v_MUX1_4844_out0[3:0];
assign v__4585_out1 = v_MUX1_4844_out0[15:12];
assign v__4586_out0 = v_MUX1_4845_out0[3:0];
assign v__4586_out1 = v_MUX1_4845_out0[15:12];
assign v__4783_out0 = { v_S_1241_out0,v_S_1247_out0 };
assign v__4798_out0 = { v_S_1465_out0,v_S_1471_out0 };
assign v_TX_INSTRUCTION_13659_out0 = v_TX_INSTRUCTION_7012_out0;
assign v_TX_INSTRUCTION_13660_out0 = v_TX_INSTRUCTION_7013_out0;
assign v_RX_INST1_12_out0 = v_RX_INSTRUCTION_2343_out0;
assign v_RX_INST0_2970_out0 = v_RX_INSTRUCTION_2344_out0;
assign v_RAMDOUT_3031_out0 = v_REGISTE_IN_4490_out0;
assign v_RAMDOUT_3032_out0 = v_REGISTE_IN_4491_out0;
assign v__4660_out0 = { v__4585_out1,v_C1_6919_out0 };
assign v__4661_out0 = { v__4586_out1,v_C1_6920_out0 };
assign v_NOTUSED_9800_out0 = v__4585_out0;
assign v_NOTUSED_9801_out0 = v__4586_out0;
assign v_CIN_9831_out0 = v_COUT_715_out0;
assign v_CIN_10055_out0 = v_COUT_939_out0;
assign v_TX_INST_10827_out0 = v_TX_INSTRUCTION_13659_out0;
assign v_TX_INST_10828_out0 = v_TX_INSTRUCTION_13660_out0;
assign v_REGISTER_INPUT_13621_out0 = v_REGISTE_IN_4490_out0;
assign v_REGISTER_INPUT_13622_out0 = v_REGISTE_IN_4491_out0;
assign v_SHIFTED_SIG_13632_out0 = v_shifted1_2666_out0;
assign v_SHIFTED_SIG_13633_out0 = v_shifted1_2667_out0;
assign v_RAMDOUT_23_out0 = v_RAMDOUT_3031_out0;
assign v_RAMDOUT_24_out0 = v_RAMDOUT_3032_out0;
assign v_REGISTER_INUP16_384_out0 = v_REGISTER_INPUT_13621_out0;
assign v_TX_INSTRUCTION1_1169_out0 = v_TX_INST_10827_out0;
assign v_TX_INSTRUCTION0_1762_out0 = v_TX_INST_10828_out0;
assign v_G1_2354_out0 = v_RX_INST1_12_out0 || v_RX_INST0_2970_out0;
assign v_RD_5912_out0 = v_CIN_9831_out0;
assign v_RD_6376_out0 = v_CIN_10055_out0;
assign v_SHIFTED_SIG_10802_out0 = v_SHIFTED_SIG_13632_out0;
assign v_SHIFTED_SIG_10803_out0 = v_SHIFTED_SIG_13633_out0;
assign v_REGISTER_INUP0_12240_out0 = v_REGISTER_INPUT_13622_out0;
assign v_MUX2_13319_out0 = v_LSR_418_out0 ? v__4660_out0 : v_MUX1_4844_out0;
assign v_MUX2_13320_out0 = v_LSR_419_out0 ? v__4661_out0 : v_MUX1_4845_out0;
assign v_MUX2_188_out0 = v_SHIFT_WHICH_OP_4459_out0 ? v_RD_SIG11_7132_out0 : v_SHIFTED_SIG_10802_out0;
assign v_MUX2_189_out0 = v_SHIFT_WHICH_OP_4460_out0 ? v_RD_SIG11_7133_out0 : v_SHIFTED_SIG_10803_out0;
assign v_TX_INSTUCTION0_228_out0 = v_TX_INSTRUCTION0_1762_out0;
assign v_RX_INST_2334_out0 = v_G1_2354_out0;
assign v_IN_2350_out0 = v_MUX2_13319_out0;
assign v_IN_2351_out0 = v_MUX2_13320_out0;
assign v_RAMDOUT_2414_out0 = v_RAMDOUT_23_out0;
assign v_RAMDOUT_2415_out0 = v_RAMDOUT_24_out0;
assign v_TX_INSTUCTION1_4859_out0 = v_TX_INSTRUCTION1_1169_out0;
assign v_MUX1_7702_out0 = v_SHIFT_WHICH_OP_4459_out0 ? v_SHIFTED_SIG_10802_out0 : v_OP2_SIG11_4827_out0;
assign v_MUX1_7703_out0 = v_SHIFT_WHICH_OP_4460_out0 ? v_SHIFTED_SIG_10803_out0 : v_OP2_SIG11_4828_out0;
assign v_G1_7767_out0 = ((v_RD_5912_out0 && !v_RM_11352_out0) || (!v_RD_5912_out0) && v_RM_11352_out0);
assign v_G1_8231_out0 = ((v_RD_6376_out0 && !v_RM_11816_out0) || (!v_RD_6376_out0) && v_RM_11816_out0);
assign v_G2_12303_out0 = v_RD_5912_out0 && v_RM_11352_out0;
assign v_G2_12767_out0 = v_RD_6376_out0 && v_RM_11816_out0;
assign v_TX_inst0_608_out0 = v_TX_INSTUCTION0_228_out0;
assign v_MUX1_1735_out0 = v_EXEC1_20_out0 ? v_RMN_13437_out0 : v_RAMDOUT_2414_out0;
assign v_MUX1_1736_out0 = v_EXEC1_21_out0 ? v_RMN_13438_out0 : v_RAMDOUT_2415_out0;
assign v_CARRY_4912_out0 = v_G2_12303_out0;
assign v_CARRY_5376_out0 = v_G2_12767_out0;
assign v_RX_INSTRUCTION_8686_out0 = v_RX_INST_2334_out0;
assign v_RD_SIG_NEW_8759_out0 = v_MUX2_188_out0;
assign v_RD_SIG_NEW_8760_out0 = v_MUX2_189_out0;
assign v_S_8913_out0 = v_G1_7767_out0;
assign v_S_9377_out0 = v_G1_8231_out0;
assign v__10536_out0 = v_IN_2350_out0[15:15];
assign v__10537_out0 = v_IN_2351_out0[15:15];
assign v_OP2_SIG_NEW_11190_out0 = v_MUX1_7702_out0;
assign v_OP2_SIG_NEW_11191_out0 = v_MUX1_7703_out0;
assign v__13291_out0 = v_IN_2350_out0[3:0];
assign v__13291_out1 = v_IN_2350_out0[15:12];
assign v__13292_out0 = v_IN_2351_out0[3:0];
assign v__13292_out1 = v_IN_2351_out0[15:12];
assign v__164_out0 = { v__13291_out1,v__10536_out0 };
assign v__165_out0 = { v__13292_out1,v__10537_out0 };
assign v_S_1242_out0 = v_S_8913_out0;
assign v_S_1466_out0 = v_S_9377_out0;
assign v_G1_4018_out0 = v_CARRY_4912_out0 || v_CARRY_4911_out0;
assign v_G1_4242_out0 = v_CARRY_5376_out0 || v_CARRY_5375_out0;
assign v_RX_INSTRUCTION_4659_out0 = v_RX_INSTRUCTION_8686_out0;
assign v_MUX5_7678_out0 = v_TX_inst0_608_out0 ? v_BYTE_COMP_10_13611_out0 : v_BYTE_COMP_11_1163_out0;
assign v_RD_SIG_NEW_10872_out0 = v_RD_SIG_NEW_8759_out0;
assign v_RD_SIG_NEW_10873_out0 = v_RD_SIG_NEW_8760_out0;
assign v_REGDIN_11041_out0 = v_MUX1_1735_out0;
assign v_REGDIN_11042_out0 = v_MUX1_1736_out0;
assign v_OP2_SIG_NEW_11218_out0 = v_OP2_SIG_NEW_11190_out0;
assign v_OP2_SIG_NEW_11219_out0 = v_OP2_SIG_NEW_11191_out0;
assign v_NOTUSED_13265_out0 = v__13291_out0;
assign v_NOTUSED_13266_out0 = v__13292_out0;
assign v_G22_13663_out0 = v_TX_inst0_608_out0 || v_TX_INSTUCTION1_4859_out0;
assign v_RD_SIG_109_out0 = v_RD_SIG_NEW_10872_out0;
assign v_RD_SIG_110_out0 = v_RD_SIG_NEW_10873_out0;
assign v_COUT_710_out0 = v_G1_4018_out0;
assign v_COUT_934_out0 = v_G1_4242_out0;
assign v__2553_out0 = { v__4783_out0,v_S_1242_out0 };
assign v__2568_out0 = { v__4798_out0,v_S_1466_out0 };
assign v_LS_REGIN_3303_out0 = v_REGDIN_11041_out0;
assign v_LS_REGIN_3304_out0 = v_REGDIN_11042_out0;
assign v_byte_comp_1_6923_out0 = v_MUX5_7678_out0;
assign v__11055_out0 = { v__164_out0,v__10536_out0 };
assign v__11056_out0 = { v__165_out0,v__10537_out0 };
assign v_TX_INST_11239_out0 = v_G22_13663_out0;
assign v_OP2_SIG_13314_out0 = v_OP2_SIG_NEW_11218_out0;
assign v_OP2_SIG_13315_out0 = v_OP2_SIG_NEW_11219_out0;
assign v_RX_INSTRUCTION_13325_out0 = v_RX_INSTRUCTION_4659_out0;
assign v__3178_out0 = { v_OP2_SIG_13314_out0,v_C4_2593_out0 };
assign v__3179_out0 = { v_OP2_SIG_13315_out0,v_C4_2594_out0 };
assign v_byte_comp_1_6872_out0 = v_byte_comp_1_6923_out0;
assign v_G4_6915_out0 = ! v_RX_INSTRUCTION_13325_out0;
assign v_G8_7103_out0 = v_RX_INSTRUCTION_13325_out0 || v_RXBYTERECEIVED_3269_out0;
assign v_CIN_9826_out0 = v_COUT_710_out0;
assign v_CIN_10050_out0 = v_COUT_934_out0;
assign v_G18_10489_out0 = ! v_RX_INSTRUCTION_13325_out0;
assign v_TX_INSTRUCTION_10501_out0 = v_TX_INST_11239_out0;
assign v__11231_out0 = { v__11055_out0,v__10536_out0 };
assign v__11232_out0 = { v__11056_out0,v__10537_out0 };
assign v__13275_out0 = { v_RD_SIG_109_out0,v_C4_2593_out0 };
assign v__13276_out0 = { v_RD_SIG_110_out0,v_C4_2594_out0 };
assign v__2791_out0 = { v__11231_out0,v__10536_out0 };
assign v__2792_out0 = { v__11232_out0,v__10537_out0 };
assign v_G3_3948_out0 = v_G4_6915_out0 && v_G1_10476_out0;
assign v_XOR2_4486_out0 = v__3178_out0 ^ v_C11_4539_out0;
assign v_XOR2_4487_out0 = v__3179_out0 ^ v_C11_4540_out0;
assign v_RD_5900_out0 = v_CIN_9826_out0;
assign v_RD_6364_out0 = v_CIN_10050_out0;
assign v_G16_7701_out0 = v_G19_3860_out0 && v_G18_10489_out0;
assign v_BYTE_COMP_1_8743_out0 = v_byte_comp_1_6872_out0;
assign v_XOR1_11246_out0 = v__13275_out0 ^ v_C5_2688_out0;
assign v_XOR1_11247_out0 = v__13276_out0 ^ v_C5_2689_out0;
assign v_TX_INSTRUCTION_13631_out0 = v_TX_INSTRUCTION_10501_out0;
assign v_OUT_460_out0 = v__2791_out0;
assign v_OUT_461_out0 = v__2792_out0;
assign {v_A5_1901_out1,v_A5_1901_out0 } = v_C7_1865_out0 + v_XOR2_4486_out0 + v_C12_1151_out0;
assign {v_A5_1902_out1,v_A5_1902_out0 } = v_C7_1866_out0 + v_XOR2_4487_out0 + v_C12_1152_out0;
assign v_TX_INSTRUCTION_6875_out0 = v_TX_INSTRUCTION_13631_out0;
assign v_G1_7755_out0 = ((v_RD_5900_out0 && !v_RM_11340_out0) || (!v_RD_5900_out0) && v_RM_11340_out0);
assign v_G1_8219_out0 = ((v_RD_6364_out0 && !v_RM_11804_out0) || (!v_RD_6364_out0) && v_RM_11804_out0);
assign v_G5_10801_out0 = v_G3_3948_out0 && v__2983_out0;
assign v_G20_11040_out0 = v_G17_1903_out0 || v_G16_7701_out0;
assign v_G7_11095_out0 = v_G6_4818_out0 && v_G3_3948_out0;
assign {v_A4_11227_out1,v_A4_11227_out0 } = v_XOR1_11246_out0 + v_C7_1865_out0 + v_C6_10317_out0;
assign {v_A4_11228_out1,v_A4_11228_out0 } = v_XOR1_11247_out0 + v_C7_1866_out0 + v_C6_10318_out0;
assign v_G2_12291_out0 = v_RD_5900_out0 && v_RM_11340_out0;
assign v_G2_12755_out0 = v_RD_6364_out0 && v_RM_11804_out0;
assign v_TX_INSTRUCTION_453_out0 = v_TX_INSTRUCTION_6875_out0;
assign v_MUX2_1181_out0 = v_G1_289_out0 ? v_A5_1901_out0 : v__3178_out0;
assign v_MUX2_1182_out0 = v_G1_290_out0 ? v_A5_1902_out0 : v__3179_out0;
assign v_MUX1_1883_out0 = v_RD_SIGN_2405_out0 ? v_A4_11227_out0 : v__13275_out0;
assign v_MUX1_1884_out0 = v_RD_SIGN_2406_out0 ? v_A4_11228_out0 : v__13276_out0;
assign v_MUX3_3041_out0 = v_ASR_10566_out0 ? v_OUT_460_out0 : v_MUX2_13319_out0;
assign v_MUX3_3042_out0 = v_ASR_10567_out0 ? v_OUT_461_out0 : v_MUX2_13320_out0;
assign v_CARRY_4900_out0 = v_G2_12291_out0;
assign v_CARRY_5364_out0 = v_G2_12755_out0;
assign v_S_8901_out0 = v_G1_7755_out0;
assign v_S_9365_out0 = v_G1_8219_out0;
assign v_NOTUSED4_10530_out0 = v_A4_11227_out1;
assign v_NOTUSED4_10531_out0 = v_A4_11228_out1;
assign v_NOTUSED1_10684_out0 = v_A5_1901_out1;
assign v_NOTUSED1_10685_out0 = v_A5_1902_out1;
assign v_G10_10694_out0 = v_G5_10801_out0 || v_G9_13655_out0;
assign v_S_1237_out0 = v_S_8901_out0;
assign v_S_1461_out0 = v_S_9365_out0;
assign v_TRANSMIT_INSTRUCTION_1713_out0 = v_TX_INSTRUCTION_453_out0;
assign v_TX_INSTRUCTION_2825_out0 = v_TX_INSTRUCTION_453_out0;
assign v_G1_4013_out0 = v_CARRY_4900_out0 || v_CARRY_4899_out0;
assign v_G1_4237_out0 = v_CARRY_5364_out0 || v_CARRY_5363_out0;
assign v__4488_out0 = v_MUX3_3041_out0[3:0];
assign v__4488_out1 = v_MUX3_3041_out0[15:12];
assign v__4489_out0 = v_MUX3_3042_out0[3:0];
assign v__4489_out1 = v_MUX3_3042_out0[15:12];
assign v__4547_out0 = { v_G7_11095_out0,v_G10_10694_out0 };
assign {v_A6_10463_out1,v_A6_10463_out0 } = v_MUX1_1883_out0 + v_MUX2_1181_out0 + v_C3_4741_out0;
assign {v_A6_10464_out1,v_A6_10464_out0 } = v_MUX1_1884_out0 + v_MUX2_1182_out0 + v_C3_4742_out0;
assign v__167_out0 = { v__4488_out1,v__4488_out0 };
assign v__168_out0 = { v__4489_out1,v__4489_out0 };
assign v_COUT_705_out0 = v_G1_4013_out0;
assign v_COUT_929_out0 = v_G1_4237_out0;
assign v_SEL1_2305_out0 = v_A6_10463_out0[15:15];
assign v_SEL1_2306_out0 = v_A6_10464_out0[15:15];
assign v_G23_2614_out0 = v_G21_10681_out0 && v_TX_INSTRUCTION_2825_out0;
assign v_transmit_INSTRUCTION_2674_out0 = v_TRANSMIT_INSTRUCTION_1713_out0;
assign v__7033_out0 = { v__2553_out0,v_S_1237_out0 };
assign v__7048_out0 = { v__2568_out0,v_S_1461_out0 };
assign v_NOTUSED_10835_out0 = v_A6_10463_out1;
assign v_NOTUSED_10836_out0 = v_A6_10464_out1;
assign v_MUX1_11061_out0 = v_RX_INSTRUCTION_13325_out0 ? v_C5_10356_out0 : v__4547_out0;
assign v_XOR3_13599_out0 = v_A6_10463_out0 ^ v_C15_1730_out0;
assign v_XOR3_13600_out0 = v_A6_10464_out0 ^ v_C15_1731_out0;
assign v_SIGN_ANS_1970_out0 = v_SEL1_2305_out0;
assign v_SIGN_ANS_1971_out0 = v_SEL1_2306_out0;
assign v_MUX4_2229_out0 = v_ROR_544_out0 ? v__167_out0 : v_MUX3_3041_out0;
assign v_MUX4_2230_out0 = v_ROR_545_out0 ? v__168_out0 : v_MUX3_3042_out0;
assign v_MUX8_2697_out0 = v_transmit_INSTRUCTION_2674_out0 ? v_C1_10259_out0 : v_FF8_11222_out0;
assign v_CIN_9825_out0 = v_COUT_705_out0;
assign v_CIN_10049_out0 = v_COUT_929_out0;
assign v_G24_10460_out0 = ! v_G23_2614_out0;
assign v_G2_10471_out0 = ! v_transmit_INSTRUCTION_2674_out0;
assign v_MUX3_10994_out0 = v_G25_4658_out0 ? v_G23_2614_out0 : v_C7_3222_out0;
assign {v_A8_11155_out1,v_A8_11155_out0 } = v_XOR3_13599_out0 + v_C13_2185_out0 + v_C14_1674_out0;
assign {v_A8_11156_out1,v_A8_11156_out0 } = v_XOR3_13600_out0 + v_C13_2186_out0 + v_C14_1675_out0;
assign v_G3_13507_out0 = v_transmit_INSTRUCTION_2674_out0 || v_SHIFHT_ENABLE_13501_out0;
assign v_TX_OVERFLOW_500_out0 = v_MUX3_10994_out0;
assign v_G10_602_out0 = v_G7_2455_out0 && v_G2_10471_out0;
assign v__1813_out0 = { v_MUX3_10994_out0,v_C4_1201_out0 };
assign v_ENABLE_2651_out0 = v_G3_13507_out0;
assign v_NOTUSED2_5794_out0 = v_A8_11155_out1;
assign v_NOTUSED2_5795_out0 = v_A8_11156_out1;
assign v_RD_5898_out0 = v_CIN_9825_out0;
assign v_RD_6362_out0 = v_CIN_10049_out0;
assign v_STARTBIT_6968_out0 = v_G2_10471_out0;
assign v_STARTBIT_6970_out0 = v_G24_10460_out0;
assign v_SIGN_ANS_8650_out0 = v_SIGN_ANS_1970_out0;
assign v_SIGN_ANS_8651_out0 = v_SIGN_ANS_1971_out0;
assign v_MUX3_8669_out0 = v_SEL1_2305_out0 ? v_A8_11155_out0 : v_A6_10463_out0;
assign v_MUX3_8670_out0 = v_SEL1_2306_out0 ? v_A8_11156_out0 : v_A6_10464_out0;
assign v_MUX5_10605_out0 = v_EN_13181_out0 ? v_MUX4_2229_out0 : v_IN_13548_out0;
assign v_MUX5_10606_out0 = v_EN_13182_out0 ? v_MUX4_2230_out0 : v_IN_13549_out0;
assign v_MUX9_166_out0 = v_G10_602_out0 ? v_2_7072_out0 : v_FF9_8805_out0;
assign v_OUT_2352_out0 = v_MUX5_10605_out0;
assign v_OUT_2353_out0 = v_MUX5_10606_out0;
assign v_SIGN_ANS_4457_out0 = v_SIGN_ANS_8650_out0;
assign v_SIGN_ANS_4458_out0 = v_SIGN_ANS_8651_out0;
assign v_G1_7753_out0 = ((v_RD_5898_out0 && !v_RM_11338_out0) || (!v_RD_5898_out0) && v_RM_11338_out0);
assign v_G1_8217_out0 = ((v_RD_6362_out0 && !v_RM_11802_out0) || (!v_RD_6362_out0) && v_RM_11802_out0);
assign v_G35_10361_out0 = v_STARTBIT_6968_out0 && v_G36_3136_out0;
assign v_G35_10363_out0 = v_STARTBIT_6970_out0 && v_G36_3138_out0;
assign v_TX_OVERFLOW_10481_out0 = v_TX_OVERFLOW_500_out0;
assign v_SEL8_10686_out0 = v_MUX3_8669_out0[11:0];
assign v_SEL8_10687_out0 = v_MUX3_8670_out0[11:0];
assign v_G2_12289_out0 = v_RD_5898_out0 && v_RM_11338_out0;
assign v_G2_12753_out0 = v_RD_6362_out0 && v_RM_11802_out0;
assign v_IN_190_out0 = v_OUT_2352_out0;
assign v_IN_191_out0 = v_OUT_2353_out0;
assign v_ENABLE_2019_out0 = v_G35_10361_out0;
assign v_ENABLE_2021_out0 = v_G35_10363_out0;
assign v_OUTSTREAM_2097_out0 = v_MUX9_166_out0;
assign v_CARRY_4898_out0 = v_G2_12289_out0;
assign v_CARRY_5362_out0 = v_G2_12753_out0;
assign v_S_8899_out0 = v_G1_7753_out0;
assign v_S_9363_out0 = v_G1_8217_out0;
assign v_SIGN_ANS_10302_out0 = v_SIGN_ANS_4457_out0;
assign v_SIGN_ANS_10303_out0 = v_SIGN_ANS_4458_out0;
assign v_TX_OVERFLOW_13294_out0 = v_TX_OVERFLOW_10481_out0;
assign v_OUT_22_out0 = v_OUTSTREAM_2097_out0;
assign v_IN_685_out0 = v_IN_190_out0;
assign v_IN_686_out0 = v_IN_191_out0;
assign v_S_1236_out0 = v_S_8899_out0;
assign v_S_1460_out0 = v_S_9363_out0;
assign v__3125_out0 = v_IN_190_out0[7:0];
assign v__3125_out1 = v_IN_190_out0[15:8];
assign v__3126_out0 = v_IN_191_out0[7:0];
assign v__3126_out1 = v_IN_191_out0[15:8];
assign v_G1_4012_out0 = v_CARRY_4898_out0 || v_CARRY_4897_out0;
assign v_G1_4236_out0 = v_CARRY_5362_out0 || v_CARRY_5361_out0;
assign v_G18_8800_out0 = !(v_ENABLE_2019_out0 || v_Q7_6889_out0);
assign v_G18_8802_out0 = !(v_ENABLE_2021_out0 || v_Q7_6891_out0);
assign v_NOTUSED2_41_out0 = v__3125_out1;
assign v_NOTUSED2_42_out0 = v__3126_out1;
assign v_COUT_704_out0 = v_G1_4012_out0;
assign v_COUT_928_out0 = v_G1_4236_out0;
assign v_BIT_OUT_2015_out0 = v_OUT_22_out0;
assign v_G21_3809_out0 = v_G18_8800_out0 || v_G22_10984_out0;
assign v_G21_3811_out0 = v_G18_8802_out0 || v_G22_10986_out0;
assign v__4709_out0 = { v_C1_13446_out0,v__3125_out0 };
assign v__4710_out0 = { v_C1_13447_out0,v__3126_out0 };
assign v__13519_out0 = { v__7033_out0,v_S_1236_out0 };
assign v__13534_out0 = { v__7048_out0,v_S_1460_out0 };
assign v_BIT_383_out0 = v_BIT_OUT_2015_out0;
assign v_CIN_9832_out0 = v_COUT_704_out0;
assign v_CIN_10056_out0 = v_COUT_928_out0;
assign v_MUX1_10443_out0 = v_LSL_1861_out0 ? v__4709_out0 : v_IN_685_out0;
assign v_MUX1_10444_out0 = v_LSL_1862_out0 ? v__4710_out0 : v_IN_686_out0;
assign v_BIT_OUT_10705_out0 = v_BIT_OUT_2015_out0;
assign v_G2_3214_out0 = ! v_BIT_383_out0;
assign v_RD_5914_out0 = v_CIN_9832_out0;
assign v_RD_6378_out0 = v_CIN_10056_out0;
assign v_STARTBIT_6969_out0 = v_BIT_383_out0;
assign v__8673_out0 = v_MUX1_10443_out0[7:0];
assign v__8673_out1 = v_MUX1_10443_out0[15:8];
assign v__8674_out0 = v_MUX1_10444_out0[7:0];
assign v__8674_out1 = v_MUX1_10444_out0[15:8];
assign v_BIT_OUT_13326_out0 = v_BIT_OUT_10705_out0;
assign v_MUX2_1180_out0 = v_G22_10620_out0 ? v_G2_3214_out0 : v_C6_1732_out0;
assign v_G1_7769_out0 = ((v_RD_5914_out0 && !v_RM_11354_out0) || (!v_RD_5914_out0) && v_RM_11354_out0);
assign v_G1_8233_out0 = ((v_RD_6378_out0 && !v_RM_11818_out0) || (!v_RD_6378_out0) && v_RM_11818_out0);
assign v_G35_10362_out0 = v_STARTBIT_6969_out0 && v_G36_3137_out0;
assign v__10504_out0 = { v__8673_out1,v_C1_13446_out0 };
assign v__10505_out0 = { v__8674_out1,v_C1_13447_out0 };
assign v_NOTUSED_10564_out0 = v__8673_out0;
assign v_NOTUSED_10565_out0 = v__8674_out0;
assign v_G2_12305_out0 = v_RD_5914_out0 && v_RM_11354_out0;
assign v_G2_12769_out0 = v_RD_6378_out0 && v_RM_11818_out0;
assign v_ENABLE_2020_out0 = v_G35_10362_out0;
assign v_MUX2_2337_out0 = v_LSR_1174_out0 ? v__10504_out0 : v_MUX1_10443_out0;
assign v_MUX2_2338_out0 = v_LSR_1175_out0 ? v__10505_out0 : v_MUX1_10444_out0;
assign v_CARRY_4914_out0 = v_G2_12305_out0;
assign v_CARRY_5378_out0 = v_G2_12769_out0;
assign v_TX_PROGRESS_8645_out0 = v_MUX2_1180_out0;
assign v_S_8915_out0 = v_G1_7769_out0;
assign v_S_9379_out0 = v_G1_8233_out0;
assign v__13337_out0 = { v_MUX2_1180_out0,v_C3_10853_out0 };
assign v_TX_IN_PROGRESS_235_out0 = v_TX_PROGRESS_8645_out0;
assign v_S_1243_out0 = v_S_8915_out0;
assign v_S_1467_out0 = v_S_9379_out0;
assign v__2425_out0 = { v__13337_out0,v__1813_out0 };
assign v_G1_4019_out0 = v_CARRY_4914_out0 || v_CARRY_4913_out0;
assign v_G1_4243_out0 = v_CARRY_5378_out0 || v_CARRY_5377_out0;
assign v_IN_5796_out0 = v_MUX2_2337_out0;
assign v_IN_5797_out0 = v_MUX2_2338_out0;
assign v_G18_8801_out0 = !(v_ENABLE_2020_out0 || v_Q7_6890_out0);
assign v_COUT_711_out0 = v_G1_4019_out0;
assign v_COUT_935_out0 = v_G1_4243_out0;
assign v__2582_out0 = v_IN_5796_out0[7:0];
assign v__2582_out1 = v_IN_5796_out0[15:8];
assign v__2583_out0 = v_IN_5797_out0[7:0];
assign v__2583_out1 = v_IN_5797_out0[15:8];
assign v__3266_out0 = v_IN_5796_out0[15:15];
assign v__3267_out0 = v_IN_5797_out0[15:15];
assign v__3312_out0 = { v__13519_out0,v_S_1243_out0 };
assign v__3327_out0 = { v__13534_out0,v_S_1467_out0 };
assign v_G21_3810_out0 = v_G18_8801_out0 || v_G22_10985_out0;
assign v__10532_out0 = { v__10376_out0,v__2425_out0 };
assign v_TX_IN_PROGRESS_13634_out0 = v_TX_IN_PROGRESS_235_out0;
assign v_NOTUSED_68_out0 = v__2582_out0;
assign v_NOTUSED_69_out0 = v__2583_out0;
assign v__7704_out0 = { v__2582_out1,v__3266_out0 };
assign v__7705_out0 = { v__2583_out1,v__3267_out0 };
assign v_CIN_9833_out0 = v_COUT_711_out0;
assign v_CIN_10057_out0 = v_COUT_935_out0;
assign v_RD_STATUS_10500_out0 = v__10532_out0;
assign v_RD_5916_out0 = v_CIN_9833_out0;
assign v_RD_6380_out0 = v_CIN_10057_out0;
assign v_STATUS_REGISTER_10359_out0 = v_RD_STATUS_10500_out0;
assign v__10806_out0 = { v__7704_out0,v__3266_out0 };
assign v__10807_out0 = { v__7705_out0,v__3267_out0 };
assign v_STATUS_REGISTER_185_out0 = v_STATUS_REGISTER_10359_out0;
assign v_G1_7771_out0 = ((v_RD_5916_out0 && !v_RM_11356_out0) || (!v_RD_5916_out0) && v_RM_11356_out0);
assign v_G1_8235_out0 = ((v_RD_6380_out0 && !v_RM_11820_out0) || (!v_RD_6380_out0) && v_RM_11820_out0);
assign v_G2_12307_out0 = v_RD_5916_out0 && v_RM_11356_out0;
assign v_G2_12771_out0 = v_RD_6380_out0 && v_RM_11820_out0;
assign v__13310_out0 = { v__10806_out0,v__3266_out0 };
assign v__13311_out0 = { v__10807_out0,v__3267_out0 };
assign v__107_out0 = { v__13310_out0,v__3266_out0 };
assign v__108_out0 = { v__13311_out0,v__3267_out0 };
assign v_CARRY_4916_out0 = v_G2_12307_out0;
assign v_CARRY_5380_out0 = v_G2_12771_out0;
assign v_S_8917_out0 = v_G1_7771_out0;
assign v_S_9381_out0 = v_G1_8235_out0;
assign v_STATUS_REGISTER_13778_out0 = v_STATUS_REGISTER_185_out0;
assign v_S_1244_out0 = v_S_8917_out0;
assign v_S_1468_out0 = v_S_9381_out0;
assign v_STATUS_REGISTER_2866_out0 = v_STATUS_REGISTER_13778_out0;
assign v_STATUS_REGISTER_2867_out0 = v_STATUS_REGISTER_13778_out0;
assign v_G1_4020_out0 = v_CARRY_4916_out0 || v_CARRY_4915_out0;
assign v_G1_4244_out0 = v_CARRY_5380_out0 || v_CARRY_5379_out0;
assign v__5851_out0 = { v__107_out0,v__3266_out0 };
assign v__5852_out0 = { v__108_out0,v__3267_out0 };
assign v__538_out0 = { v__5851_out0,v__3266_out0 };
assign v__539_out0 = { v__5852_out0,v__3267_out0 };
assign v_COUT_712_out0 = v_G1_4020_out0;
assign v_COUT_936_out0 = v_G1_4244_out0;
assign v_STATUS_REGISTER_5858_out0 = v_STATUS_REGISTER_2866_out0;
assign v_STATUS_REGISTER_5859_out0 = v_STATUS_REGISTER_2867_out0;
assign v__7148_out0 = { v__3312_out0,v_S_1244_out0 };
assign v__7163_out0 = { v__3327_out0,v_S_1468_out0 };
assign v__2223_out0 = { v__538_out0,v__3266_out0 };
assign v__2224_out0 = { v__539_out0,v__3267_out0 };
assign v_MUX4_4579_out0 = v_STAT_INSTRUCTION_2855_out0 ? v_STATUS_REGISTER_5858_out0 : v_RAM_OUT_11214_out0;
assign v_MUX4_4580_out0 = v_STAT_INSTRUCTION_2856_out0 ? v_STATUS_REGISTER_5859_out0 : v_RAM_OUT_11215_out0;
assign v_CIN_9835_out0 = v_COUT_712_out0;
assign v_CIN_10059_out0 = v_COUT_936_out0;
assign v_DFQDF_3025_out0 = v_MUX4_4579_out0;
assign v_DFQDF_3026_out0 = v_MUX4_4580_out0;
assign v_RD_5920_out0 = v_CIN_9835_out0;
assign v_RD_6384_out0 = v_CIN_10059_out0;
assign v__7124_out0 = { v__2223_out0,v__3266_out0 };
assign v__7125_out0 = { v__2224_out0,v__3267_out0 };
assign v_OUT_2857_out0 = v__7124_out0;
assign v_OUT_2858_out0 = v__7125_out0;
assign v_G1_7775_out0 = ((v_RD_5920_out0 && !v_RM_11360_out0) || (!v_RD_5920_out0) && v_RM_11360_out0);
assign v_G1_8239_out0 = ((v_RD_6384_out0 && !v_RM_11824_out0) || (!v_RD_6384_out0) && v_RM_11824_out0);
assign v_G2_12311_out0 = v_RD_5920_out0 && v_RM_11360_out0;
assign v_G2_12775_out0 = v_RD_6384_out0 && v_RM_11824_out0;
assign v_CARRY_4920_out0 = v_G2_12311_out0;
assign v_CARRY_5384_out0 = v_G2_12775_out0;
assign v_MUX3_6864_out0 = v_ASR_10366_out0 ? v_OUT_2857_out0 : v_MUX2_2337_out0;
assign v_MUX3_6865_out0 = v_ASR_10367_out0 ? v_OUT_2858_out0 : v_MUX2_2338_out0;
assign v_S_8921_out0 = v_G1_7775_out0;
assign v_S_9385_out0 = v_G1_8239_out0;
assign v_S_1246_out0 = v_S_8921_out0;
assign v_S_1470_out0 = v_S_9385_out0;
assign v_G1_4022_out0 = v_CARRY_4920_out0 || v_CARRY_4919_out0;
assign v_G1_4246_out0 = v_CARRY_5384_out0 || v_CARRY_5383_out0;
assign v__11132_out0 = v_MUX3_6864_out0[7:0];
assign v__11132_out1 = v_MUX3_6864_out0[15:8];
assign v__11133_out0 = v_MUX3_6865_out0[7:0];
assign v__11133_out1 = v_MUX3_6865_out0[15:8];
assign v_COUT_714_out0 = v_G1_4022_out0;
assign v_COUT_938_out0 = v_G1_4246_out0;
assign v__4750_out0 = { v__7148_out0,v_S_1246_out0 };
assign v__4765_out0 = { v__7163_out0,v_S_1470_out0 };
assign v__6870_out0 = { v__11132_out1,v__11132_out0 };
assign v__6871_out0 = { v__11133_out1,v__11133_out0 };
assign v_CIN_9828_out0 = v_COUT_714_out0;
assign v_CIN_10052_out0 = v_COUT_938_out0;
assign v_MUX4_13498_out0 = v_ROR_282_out0 ? v__6870_out0 : v_MUX3_6864_out0;
assign v_MUX4_13499_out0 = v_ROR_283_out0 ? v__6871_out0 : v_MUX3_6865_out0;
assign v_MUX5_3305_out0 = v_EN_2445_out0 ? v_MUX4_13498_out0 : v_IN_685_out0;
assign v_MUX5_3306_out0 = v_EN_2446_out0 ? v_MUX4_13499_out0 : v_IN_686_out0;
assign v_RD_5906_out0 = v_CIN_9828_out0;
assign v_RD_6370_out0 = v_CIN_10052_out0;
assign v_G1_7761_out0 = ((v_RD_5906_out0 && !v_RM_11346_out0) || (!v_RD_5906_out0) && v_RM_11346_out0);
assign v_G1_8225_out0 = ((v_RD_6370_out0 && !v_RM_11810_out0) || (!v_RD_6370_out0) && v_RM_11810_out0);
assign v_OUT_10264_out0 = v_MUX5_3305_out0;
assign v_OUT_10265_out0 = v_MUX5_3306_out0;
assign v_G2_12297_out0 = v_RD_5906_out0 && v_RM_11346_out0;
assign v_G2_12761_out0 = v_RD_6370_out0 && v_RM_11810_out0;
assign v_OP2_2862_out0 = v_OUT_10264_out0;
assign v_OP2_2863_out0 = v_OUT_10265_out0;
assign v_CARRY_4906_out0 = v_G2_12297_out0;
assign v_CARRY_5370_out0 = v_G2_12761_out0;
assign v_S_8907_out0 = v_G1_7761_out0;
assign v_S_9371_out0 = v_G1_8225_out0;
assign v_S_1239_out0 = v_S_8907_out0;
assign v_S_1463_out0 = v_S_9371_out0;
assign v_G1_4015_out0 = v_CARRY_4906_out0 || v_CARRY_4905_out0;
assign v_G1_4239_out0 = v_CARRY_5370_out0 || v_CARRY_5369_out0;
assign v_OP2_11153_out0 = v_OP2_2862_out0;
assign v_OP2_11154_out0 = v_OP2_2863_out0;
assign v_COUT_707_out0 = v_G1_4015_out0;
assign v_COUT_931_out0 = v_G1_4239_out0;
assign v_OP2_3940_out0 = v_OP2_11153_out0;
assign v_OP2_3941_out0 = v_OP2_11154_out0;
assign v__6927_out0 = { v__4750_out0,v_S_1239_out0 };
assign v__6942_out0 = { v__4765_out0,v_S_1463_out0 };
assign v_OP2_2322_out0 = v_OP2_3940_out0;
assign v_OP2_2323_out0 = v_OP2_3941_out0;
assign v_CIN_9829_out0 = v_COUT_707_out0;
assign v_CIN_10053_out0 = v_COUT_931_out0;
assign v_RD_5908_out0 = v_CIN_9829_out0;
assign v_RD_6372_out0 = v_CIN_10053_out0;
assign v_OP2_10751_out0 = v_OP2_2322_out0;
assign v_OP2_10752_out0 = v_OP2_2323_out0;
assign v_MUX5_2595_out0 = v_MOV_196_out0 ? v_OP2_10751_out0 : v_OP1_2060_out0;
assign v_MUX5_2596_out0 = v_MOV_197_out0 ? v_OP2_10752_out0 : v_OP1_2061_out0;
assign v_B_3350_out0 = v_OP2_10751_out0;
assign v_B_3352_out0 = v_OP2_10752_out0;
assign v_G1_7763_out0 = ((v_RD_5908_out0 && !v_RM_11348_out0) || (!v_RD_5908_out0) && v_RM_11348_out0);
assign v_G1_8227_out0 = ((v_RD_6372_out0 && !v_RM_11812_out0) || (!v_RD_6372_out0) && v_RM_11812_out0);
assign v_A_11250_out0 = v_OP2_10751_out0;
assign v_A_11252_out0 = v_OP2_10752_out0;
assign v_G2_12299_out0 = v_RD_5908_out0 && v_RM_11348_out0;
assign v_G2_12763_out0 = v_RD_6372_out0 && v_RM_11812_out0;
assign v__77_out0 = v_A_11250_out0[3:3];
assign v__79_out0 = v_A_11252_out0[3:3];
assign v__192_out0 = v_A_11250_out0[15:15];
assign v__194_out0 = v_A_11252_out0[15:15];
assign v__198_out0 = v_B_3350_out0[7:7];
assign v__199_out0 = v_B_3352_out0[7:7];
assign v__321_out0 = v_A_11250_out0[0:0];
assign v__323_out0 = v_A_11252_out0[0:0];
assign v__329_out0 = v_A_11250_out0[9:9];
assign v__331_out0 = v_A_11252_out0[9:9];
assign v__1722_out0 = v_B_3350_out0[5:5];
assign v__1723_out0 = v_B_3352_out0[5:5];
assign v__1904_out0 = v_B_3350_out0[9:9];
assign v__1905_out0 = v_B_3352_out0[9:9];
assign v__2093_out0 = v_A_11250_out0[13:13];
assign v__2095_out0 = v_A_11252_out0[13:13];
assign v__2418_out0 = v_A_11250_out0[6:6];
assign v__2420_out0 = v_A_11252_out0[6:6];
assign v__2462_out0 = v_B_3350_out0[2:2];
assign v__2463_out0 = v_B_3352_out0[2:2];
assign v__2943_out0 = v_B_3350_out0[10:10];
assign v__2944_out0 = v_B_3352_out0[10:10];
assign v__3119_out0 = v_A_11250_out0[14:14];
assign v__3121_out0 = v_A_11252_out0[14:14];
assign v__3237_out0 = v_B_3350_out0[11:11];
assign v__3238_out0 = v_B_3352_out0[11:11];
assign v__3282_out0 = v_A_11250_out0[2:2];
assign v__3284_out0 = v_A_11252_out0[2:2];
assign v__4610_out0 = v_B_3350_out0[3:3];
assign v__4611_out0 = v_B_3352_out0[3:3];
assign v__4812_out0 = v_B_3350_out0[4:4];
assign v__4813_out0 = v_B_3352_out0[4:4];
assign v__4814_out0 = v_B_3350_out0[14:14];
assign v__4815_out0 = v_B_3352_out0[14:14];
assign v__4833_out0 = v_B_3350_out0[6:6];
assign v__4834_out0 = v_B_3352_out0[6:6];
assign v_CARRY_4908_out0 = v_G2_12299_out0;
assign v_CARRY_5372_out0 = v_G2_12763_out0;
assign v__7070_out0 = v_B_3350_out0[0:0];
assign v__7071_out0 = v_B_3352_out0[0:0];
assign v__8748_out0 = v_A_11250_out0[8:8];
assign v__8750_out0 = v_A_11252_out0[8:8];
assign v__8827_out0 = v_A_11250_out0[7:7];
assign v__8829_out0 = v_A_11252_out0[7:7];
assign v__8831_out0 = v_B_3350_out0[15:15];
assign v__8832_out0 = v_B_3352_out0[15:15];
assign v_S_8909_out0 = v_G1_7763_out0;
assign v_S_9373_out0 = v_G1_8227_out0;
assign v__10377_out0 = v_A_11250_out0[5:5];
assign v__10379_out0 = v_A_11252_out0[5:5];
assign v__10385_out0 = v_A_11250_out0[1:1];
assign v__10387_out0 = v_A_11252_out0[1:1];
assign v__10538_out0 = v_B_3350_out0[13:13];
assign v__10539_out0 = v_B_3352_out0[13:13];
assign v__10695_out0 = v_A_11250_out0[4:4];
assign v__10697_out0 = v_A_11252_out0[4:4];
assign v__10777_out0 = v_A_11250_out0[12:12];
assign v__10779_out0 = v_A_11252_out0[12:12];
assign v__10862_out0 = v_A_11250_out0[10:10];
assign v__10864_out0 = v_A_11252_out0[10:10];
assign v__11212_out0 = v_B_3350_out0[12:12];
assign v__11213_out0 = v_B_3352_out0[12:12];
assign v__13251_out0 = v_B_3350_out0[1:1];
assign v__13252_out0 = v_B_3352_out0[1:1];
assign v__13392_out0 = v_B_3350_out0[8:8];
assign v__13393_out0 = v_B_3352_out0[8:8];
assign v__13552_out0 = v_A_11250_out0[11:11];
assign v__13554_out0 = v_A_11252_out0[11:11];
assign v_G3_206_out0 = ((v__3282_out0 && !v_SUB_4616_out0) || (!v__3282_out0) && v_SUB_4616_out0);
assign v_G3_208_out0 = ((v__3284_out0 && !v_SUB_4618_out0) || (!v__3284_out0) && v_SUB_4618_out0);
assign v_G8_549_out0 = v__13385_out0 && v__198_out0;
assign v_G8_551_out0 = v__13387_out0 && v__199_out0;
assign v_G14_616_out0 = v__4712_out0 && v__10538_out0;
assign v_G14_618_out0 = v__4714_out0 && v__10539_out0;
assign v_G13_643_out0 = v__2876_out0 && v__11212_out0;
assign v_G13_645_out0 = v__2878_out0 && v__11213_out0;
assign v_G8_1215_out0 = ((v__8827_out0 && !v_SUB_4616_out0) || (!v__8827_out0) && v_SUB_4616_out0);
assign v_G8_1217_out0 = ((v__8829_out0 && !v_SUB_4618_out0) || (!v__8829_out0) && v_SUB_4618_out0);
assign v_S_1240_out0 = v_S_8909_out0;
assign v_S_1464_out0 = v_S_9373_out0;
assign v_G2_1810_out0 = v__13513_out0 && v__13251_out0;
assign v_G2_1812_out0 = v__13515_out0 && v__13252_out0;
assign v_G15_1814_out0 = ((v__3119_out0 && !v_SUB_4616_out0) || (!v__3119_out0) && v_SUB_4616_out0);
assign v_G15_1816_out0 = ((v__3121_out0 && !v_SUB_4618_out0) || (!v__3121_out0) && v_SUB_4618_out0);
assign v_G1_1880_out0 = v__1894_out0 && v__7070_out0;
assign v_G1_1882_out0 = v__1896_out0 && v__7071_out0;
assign v_G10_2641_out0 = v__13628_out0 && v__1904_out0;
assign v_G10_2643_out0 = v__13630_out0 && v__1905_out0;
assign v_G4_2768_out0 = v__2880_out0 && v__4610_out0;
assign v_G4_2770_out0 = v__2882_out0 && v__4611_out0;
assign v_G7_2779_out0 = ((v__2418_out0 && !v_SUB_4616_out0) || (!v__2418_out0) && v_SUB_4616_out0);
assign v_G7_2781_out0 = ((v__2420_out0 && !v_SUB_4618_out0) || (!v__2420_out0) && v_SUB_4618_out0);
assign v_G5_2784_out0 = v__1_out0 && v__4812_out0;
assign v_G5_2786_out0 = v__3_out0 && v__4813_out0;
assign v_G9_2896_out0 = v__3248_out0 && v__13392_out0;
assign v_G9_2898_out0 = v__3250_out0 && v__13393_out0;
assign v_G11_2938_out0 = v__4598_out0 && v__2943_out0;
assign v_G11_2940_out0 = v__4600_out0 && v__2944_out0;
assign v_G12_3345_out0 = ((v__13552_out0 && !v_SUB_4616_out0) || (!v__13552_out0) && v_SUB_4616_out0);
assign v_G12_3347_out0 = ((v__13554_out0 && !v_SUB_4618_out0) || (!v__13554_out0) && v_SUB_4618_out0);
assign v_G1_4016_out0 = v_CARRY_4908_out0 || v_CARRY_4907_out0;
assign v_G1_4240_out0 = v_CARRY_5372_out0 || v_CARRY_5371_out0;
assign v_G14_4533_out0 = ((v__2093_out0 && !v_SUB_4616_out0) || (!v__2093_out0) && v_SUB_4616_out0);
assign v_G14_4535_out0 = ((v__2095_out0 && !v_SUB_4618_out0) || (!v__2095_out0) && v_SUB_4618_out0);
assign v_G15_4655_out0 = v__8849_out0 && v__4814_out0;
assign v_G15_4657_out0 = v__8851_out0 && v__4815_out0;
assign v_G13_4705_out0 = ((v__10777_out0 && !v_SUB_4616_out0) || (!v__10777_out0) && v_SUB_4616_out0);
assign v_G13_4707_out0 = ((v__10779_out0 && !v_SUB_4618_out0) || (!v__10779_out0) && v_SUB_4618_out0);
assign v_G2_7025_out0 = ((v__10385_out0 && !v_SUB_4616_out0) || (!v__10385_out0) && v_SUB_4616_out0);
assign v_G2_7027_out0 = ((v__10387_out0 && !v_SUB_4618_out0) || (!v__10387_out0) && v_SUB_4618_out0);
assign v_G3_7088_out0 = v__2151_out0 && v__2462_out0;
assign v_G3_7090_out0 = v__2153_out0 && v__2463_out0;
assign v_G7_8656_out0 = v__11150_out0 && v__4833_out0;
assign v_G7_8658_out0 = v__11152_out0 && v__4834_out0;
assign v_G6_8835_out0 = v__1693_out0 && v__1722_out0;
assign v_G6_8837_out0 = v__1695_out0 && v__1723_out0;
assign v_G5_10568_out0 = ((v__10695_out0 && !v_SUB_4616_out0) || (!v__10695_out0) && v_SUB_4616_out0);
assign v_G5_10570_out0 = ((v__10697_out0 && !v_SUB_4618_out0) || (!v__10697_out0) && v_SUB_4618_out0);
assign v_G12_10689_out0 = v__1748_out0 && v__3237_out0;
assign v_G12_10691_out0 = v__1750_out0 && v__3238_out0;
assign v_G16_10907_out0 = v__2761_out0 && v__8831_out0;
assign v_G16_10909_out0 = v__2763_out0 && v__8832_out0;
assign v_G4_10997_out0 = ((v__77_out0 && !v_SUB_4616_out0) || (!v__77_out0) && v_SUB_4616_out0);
assign v_G4_10999_out0 = ((v__79_out0 && !v_SUB_4618_out0) || (!v__79_out0) && v_SUB_4618_out0);
assign v_G16_11034_out0 = ((v__192_out0 && !v_SUB_4616_out0) || (!v__192_out0) && v_SUB_4616_out0);
assign v_G16_11036_out0 = ((v__194_out0 && !v_SUB_4618_out0) || (!v__194_out0) && v_SUB_4618_out0);
assign v_G10_13215_out0 = ((v__329_out0 && !v_SUB_4616_out0) || (!v__329_out0) && v_SUB_4616_out0);
assign v_G10_13217_out0 = ((v__331_out0 && !v_SUB_4618_out0) || (!v__331_out0) && v_SUB_4618_out0);
assign v_G9_13285_out0 = ((v__8748_out0 && !v_SUB_4616_out0) || (!v__8748_out0) && v_SUB_4616_out0);
assign v_G9_13287_out0 = ((v__8750_out0 && !v_SUB_4618_out0) || (!v__8750_out0) && v_SUB_4618_out0);
assign v_G11_13342_out0 = ((v__10862_out0 && !v_SUB_4616_out0) || (!v__10862_out0) && v_SUB_4616_out0);
assign v_G11_13344_out0 = ((v__10864_out0 && !v_SUB_4618_out0) || (!v__10864_out0) && v_SUB_4618_out0);
assign v_G6_13637_out0 = ((v__10377_out0 && !v_SUB_4616_out0) || (!v__10377_out0) && v_SUB_4616_out0);
assign v_G6_13639_out0 = ((v__10379_out0 && !v_SUB_4618_out0) || (!v__10379_out0) && v_SUB_4618_out0);
assign v_G1_13757_out0 = ((v__321_out0 && !v_SUB_4616_out0) || (!v__321_out0) && v_SUB_4616_out0);
assign v_G1_13759_out0 = ((v__323_out0 && !v_SUB_4618_out0) || (!v__323_out0) && v_SUB_4618_out0);
assign v__387_out0 = { v_G5_2784_out0,v_G6_8835_out0 };
assign v__389_out0 = { v_G5_2786_out0,v_G6_8837_out0 };
assign v__400_out0 = { v_G9_2896_out0,v_G10_2641_out0 };
assign v__402_out0 = { v_G9_2898_out0,v_G10_2643_out0 };
assign v_COUT_708_out0 = v_G1_4016_out0;
assign v_COUT_932_out0 = v_G1_4240_out0;
assign v__1951_out0 = { v_G1_13757_out0,v_G2_7025_out0 };
assign v__1953_out0 = { v_G1_13759_out0,v_G2_7027_out0 };
assign v__2946_out0 = { v_G15_4655_out0,v_G16_10907_out0 };
assign v__2948_out0 = { v_G15_4657_out0,v_G16_10909_out0 };
assign v__3216_out0 = { v_G1_1880_out0,v_G2_1810_out0 };
assign v__3218_out0 = { v_G1_1882_out0,v_G2_1812_out0 };
assign v__3279_out0 = { v_G3_7088_out0,v_G4_2768_out0 };
assign v__3281_out0 = { v_G3_7090_out0,v_G4_2770_out0 };
assign v__5803_out0 = { v__6927_out0,v_S_1240_out0 };
assign v__5818_out0 = { v__6942_out0,v_S_1464_out0 };
assign v__7136_out0 = { v_G13_643_out0,v_G14_616_out0 };
assign v__7138_out0 = { v_G13_645_out0,v_G14_618_out0 };
assign v__13262_out0 = { v_G11_2938_out0,v_G12_10689_out0 };
assign v__13264_out0 = { v_G11_2940_out0,v_G12_10691_out0 };
assign v__13771_out0 = { v_G7_8656_out0,v_G8_549_out0 };
assign v__13773_out0 = { v_G7_8658_out0,v_G8_551_out0 };
assign v__114_out0 = { v__387_out0,v__13771_out0 };
assign v__116_out0 = { v__389_out0,v__13773_out0 };
assign v__450_out0 = { v__7136_out0,v__2946_out0 };
assign v__452_out0 = { v__7138_out0,v__2948_out0 };
assign v__2346_out0 = { v__400_out0,v__13262_out0 };
assign v__2348_out0 = { v__402_out0,v__13264_out0 };
assign v__9804_out0 = { v__1951_out0,v_G3_206_out0 };
assign v__9806_out0 = { v__1953_out0,v_G3_208_out0 };
assign v_CIN_9834_out0 = v_COUT_708_out0;
assign v_CIN_10058_out0 = v_COUT_932_out0;
assign v__10373_out0 = { v__3216_out0,v__3279_out0 };
assign v__10375_out0 = { v__3218_out0,v__3281_out0 };
assign v__2685_out0 = { v__10373_out0,v__114_out0 };
assign v__2687_out0 = { v__10375_out0,v__116_out0 };
assign v__4450_out0 = { v__2346_out0,v__450_out0 };
assign v__4452_out0 = { v__2348_out0,v__452_out0 };
assign v_RD_5918_out0 = v_CIN_9834_out0;
assign v_RD_6382_out0 = v_CIN_10058_out0;
assign v__8687_out0 = { v__9804_out0,v_G4_10997_out0 };
assign v__8689_out0 = { v__9806_out0,v_G4_10999_out0 };
assign v__1868_out0 = { v__2685_out0,v__4450_out0 };
assign v__1870_out0 = { v__2687_out0,v__4452_out0 };
assign v__3251_out0 = { v__8687_out0,v_G5_10568_out0 };
assign v__3253_out0 = { v__8689_out0,v_G5_10570_out0 };
assign v_G1_7773_out0 = ((v_RD_5918_out0 && !v_RM_11358_out0) || (!v_RD_5918_out0) && v_RM_11358_out0);
assign v_G1_8237_out0 = ((v_RD_6382_out0 && !v_RM_11822_out0) || (!v_RD_6382_out0) && v_RM_11822_out0);
assign v_G2_12309_out0 = v_RD_5918_out0 && v_RM_11358_out0;
assign v_G2_12773_out0 = v_RD_6382_out0 && v_RM_11822_out0;
assign v_ANDOUT_631_out0 = v__1868_out0;
assign v_ANDOUT_633_out0 = v__1870_out0;
assign v_CARRY_4918_out0 = v_G2_12309_out0;
assign v_CARRY_5382_out0 = v_G2_12773_out0;
assign v_S_8919_out0 = v_G1_7773_out0;
assign v_S_9383_out0 = v_G1_8237_out0;
assign v__10298_out0 = { v__3251_out0,v_G6_13637_out0 };
assign v__10300_out0 = { v__3253_out0,v_G6_13639_out0 };
assign v__119_out0 = { v__10298_out0,v_G7_2779_out0 };
assign v__121_out0 = { v__10300_out0,v_G7_2781_out0 };
assign v_S_1245_out0 = v_S_8919_out0;
assign v_S_1469_out0 = v_S_9383_out0;
assign v_G1_4021_out0 = v_CARRY_4918_out0 || v_CARRY_4917_out0;
assign v_G1_4245_out0 = v_CARRY_5382_out0 || v_CARRY_5381_out0;
assign v_COUT_713_out0 = v_G1_4021_out0;
assign v_COUT_937_out0 = v_G1_4245_out0;
assign v__2027_out0 = { v__5803_out0,v_S_1245_out0 };
assign v__2042_out0 = { v__5818_out0,v_S_1469_out0 };
assign v__13790_out0 = { v__119_out0,v_G8_1215_out0 };
assign v__13792_out0 = { v__121_out0,v_G8_1217_out0 };
assign v__464_out0 = { v__13790_out0,v_G9_13285_out0 };
assign v__466_out0 = { v__13792_out0,v_G9_13287_out0 };
assign v_CIN_9823_out0 = v_COUT_713_out0;
assign v_CIN_10047_out0 = v_COUT_937_out0;
assign v__422_out0 = { v__464_out0,v_G10_13215_out0 };
assign v__424_out0 = { v__466_out0,v_G10_13217_out0 };
assign v_RD_5894_out0 = v_CIN_9823_out0;
assign v_RD_6358_out0 = v_CIN_10047_out0;
assign v__2834_out0 = { v__422_out0,v_G11_13342_out0 };
assign v__2836_out0 = { v__424_out0,v_G11_13344_out0 };
assign v_G1_7749_out0 = ((v_RD_5894_out0 && !v_RM_11334_out0) || (!v_RD_5894_out0) && v_RM_11334_out0);
assign v_G1_8213_out0 = ((v_RD_6358_out0 && !v_RM_11798_out0) || (!v_RD_6358_out0) && v_RM_11798_out0);
assign v_G2_12285_out0 = v_RD_5894_out0 && v_RM_11334_out0;
assign v_G2_12749_out0 = v_RD_6358_out0 && v_RM_11798_out0;
assign v_CARRY_4894_out0 = v_G2_12285_out0;
assign v_CARRY_5358_out0 = v_G2_12749_out0;
assign v_S_8895_out0 = v_G1_7749_out0;
assign v_S_9359_out0 = v_G1_8213_out0;
assign v__11137_out0 = { v__2834_out0,v_G12_3345_out0 };
assign v__11139_out0 = { v__2836_out0,v_G12_3347_out0 };
assign v_S_1234_out0 = v_S_8895_out0;
assign v_S_1458_out0 = v_S_9359_out0;
assign v__3192_out0 = { v__11137_out0,v_G13_4705_out0 };
assign v__3194_out0 = { v__11139_out0,v_G13_4707_out0 };
assign v_G1_4010_out0 = v_CARRY_4894_out0 || v_CARRY_4893_out0;
assign v_G1_4234_out0 = v_CARRY_5358_out0 || v_CARRY_5357_out0;
assign v__173_out0 = { v__3192_out0,v_G14_4533_out0 };
assign v__175_out0 = { v__3194_out0,v_G14_4535_out0 };
assign v_COUT_702_out0 = v_G1_4010_out0;
assign v_COUT_926_out0 = v_G1_4234_out0;
assign v__2794_out0 = { v__2027_out0,v_S_1234_out0 };
assign v__2809_out0 = { v__2042_out0,v_S_1458_out0 };
assign v_CIN_9827_out0 = v_COUT_702_out0;
assign v_CIN_10051_out0 = v_COUT_926_out0;
assign v__10455_out0 = { v__173_out0,v_G15_1814_out0 };
assign v__10457_out0 = { v__175_out0,v_G15_1816_out0 };
assign v__1211_out0 = { v__10455_out0,v_G16_11034_out0 };
assign v__1213_out0 = { v__10457_out0,v_G16_11036_out0 };
assign v_RD_5902_out0 = v_CIN_9827_out0;
assign v_RD_6366_out0 = v_CIN_10051_out0;
assign v_G1_7757_out0 = ((v_RD_5902_out0 && !v_RM_11342_out0) || (!v_RD_5902_out0) && v_RM_11342_out0);
assign v_G1_8221_out0 = ((v_RD_6366_out0 && !v_RM_11806_out0) || (!v_RD_6366_out0) && v_RM_11806_out0);
assign v_ADDER_IN_8744_out0 = v__1211_out0;
assign v_ADDER_IN_8746_out0 = v__1213_out0;
assign v_G2_12293_out0 = v_RD_5902_out0 && v_RM_11342_out0;
assign v_G2_12757_out0 = v_RD_6366_out0 && v_RM_11806_out0;
assign {v_A1_3855_out1,v_A1_3855_out0 } = v_OP1_2060_out0 + v_ADDER_IN_8744_out0 + v_G10_130_out0;
assign {v_A1_3856_out1,v_A1_3856_out0 } = v_OP1_2061_out0 + v_ADDER_IN_8746_out0 + v_G10_131_out0;
assign v_CARRY_4902_out0 = v_G2_12293_out0;
assign v_CARRY_5366_out0 = v_G2_12757_out0;
assign v_S_8903_out0 = v_G1_7757_out0;
assign v_S_9367_out0 = v_G1_8221_out0;
assign v_S_1238_out0 = v_S_8903_out0;
assign v_S_1462_out0 = v_S_9367_out0;
assign v_COUT_3895_out0 = v_A1_3855_out1;
assign v_COUT_3896_out0 = v_A1_3856_out1;
assign v_G1_4014_out0 = v_CARRY_4902_out0 || v_CARRY_4901_out0;
assign v_G1_4238_out0 = v_CARRY_5366_out0 || v_CARRY_5365_out0;
assign v_SUM1_13213_out0 = v_A1_3855_out0;
assign v_SUM1_13214_out0 = v_A1_3856_out0;
assign v_COUT_706_out0 = v_G1_4014_out0;
assign v_COUT_930_out0 = v_G1_4238_out0;
assign v__1826_out0 = { v__2794_out0,v_S_1238_out0 };
assign v__1841_out0 = { v__2809_out0,v_S_1462_out0 };
assign v_MUX3_2058_out0 = v_G7_169_out0 ? v_SUM1_13213_out0 : v_MUX5_2595_out0;
assign v_MUX3_2059_out0 = v_G7_170_out0 ? v_SUM1_13214_out0 : v_MUX5_2596_out0;
assign v_MUX2_1199_out0 = v_G9_411_out0 ? v_ANDOUT_631_out0 : v_MUX3_2058_out0;
assign v_MUX2_1200_out0 = v_G9_412_out0 ? v_ANDOUT_633_out0 : v_MUX3_2059_out0;
assign v_CIN_9824_out0 = v_COUT_706_out0;
assign v_CIN_10048_out0 = v_COUT_930_out0;
assign v_RD_5896_out0 = v_CIN_9824_out0;
assign v_RD_6360_out0 = v_CIN_10048_out0;
assign v_ALUOUT_10528_out0 = v_MUX2_1199_out0;
assign v_ALUOUT_10529_out0 = v_MUX2_1200_out0;
assign v_G1_7751_out0 = ((v_RD_5896_out0 && !v_RM_11336_out0) || (!v_RD_5896_out0) && v_RM_11336_out0);
assign v_G1_8215_out0 = ((v_RD_6360_out0 && !v_RM_11800_out0) || (!v_RD_6360_out0) && v_RM_11800_out0);
assign v_ALUOUT_8856_out0 = v_ALUOUT_10528_out0;
assign v_ALUOUT_8857_out0 = v_ALUOUT_10529_out0;
assign v_G2_12287_out0 = v_RD_5896_out0 && v_RM_11336_out0;
assign v_G2_12751_out0 = v_RD_6360_out0 && v_RM_11800_out0;
assign v_ALUOUT_4607_out0 = v_ALUOUT_8856_out0;
assign v_ALUOUT_4608_out0 = v_ALUOUT_8857_out0;
assign v_CARRY_4896_out0 = v_G2_12287_out0;
assign v_CARRY_5360_out0 = v_G2_12751_out0;
assign v_S_8897_out0 = v_G1_7751_out0;
assign v_S_9361_out0 = v_G1_8215_out0;
assign v_S_1235_out0 = v_S_8897_out0;
assign v_S_1459_out0 = v_S_9361_out0;
assign v_G1_4011_out0 = v_CARRY_4896_out0 || v_CARRY_4895_out0;
assign v_G1_4235_out0 = v_CARRY_5360_out0 || v_CARRY_5359_out0;
assign v_ALUOUT_11053_out0 = v_ALUOUT_4607_out0;
assign v_ALUOUT_11054_out0 = v_ALUOUT_4608_out0;
assign v_COUT_703_out0 = v_G1_4011_out0;
assign v_COUT_927_out0 = v_G1_4235_out0;
assign v_ALUOUT_4494_out0 = v_ALUOUT_11053_out0;
assign v_ALUOUT_4495_out0 = v_ALUOUT_11054_out0;
assign v__4550_out0 = { v__1826_out0,v_S_1235_out0 };
assign v__4565_out0 = { v__1841_out0,v_S_1459_out0 };
assign v_EQ3_11044_out0 = v_ALUOUT_4494_out0 == 16'h0;
assign v_EQ3_11045_out0 = v_ALUOUT_4495_out0 == 16'h0;
assign v__11294_out0 = v_ALUOUT_4494_out0[14:0];
assign v__11294_out1 = v_ALUOUT_4494_out0[15:1];
assign v__11295_out0 = v_ALUOUT_4495_out0[14:0];
assign v__11295_out1 = v_ALUOUT_4495_out0[15:1];
assign v_RM_11344_out0 = v_COUT_703_out0;
assign v_RM_11808_out0 = v_COUT_927_out0;
assign v_EQ_100_out0 = v_EQ3_11044_out0;
assign v_EQ_101_out0 = v_EQ3_11045_out0;
assign v_REST_162_out0 = v__11294_out0;
assign v_REST_163_out0 = v__11295_out0;
assign v_MI_2612_out0 = v__11294_out1;
assign v_MI_2613_out0 = v__11295_out1;
assign v_G1_7759_out0 = ((v_RD_5904_out0 && !v_RM_11344_out0) || (!v_RD_5904_out0) && v_RM_11344_out0);
assign v_G1_8223_out0 = ((v_RD_6368_out0 && !v_RM_11808_out0) || (!v_RD_6368_out0) && v_RM_11808_out0);
assign v_G2_12295_out0 = v_RD_5904_out0 && v_RM_11344_out0;
assign v_G2_12759_out0 = v_RD_6368_out0 && v_RM_11808_out0;
assign v_MI_560_out0 = v_MI_2612_out0;
assign v_MI_561_out0 = v_MI_2613_out0;
assign v_EQ_2591_out0 = v_EQ_100_out0;
assign v_EQ_2592_out0 = v_EQ_101_out0;
assign v_CARRY_4904_out0 = v_G2_12295_out0;
assign v_CARRY_5368_out0 = v_G2_12759_out0;
assign v_S_8905_out0 = v_G1_7759_out0;
assign v_S_9369_out0 = v_G1_8223_out0;
assign v_EQ_3821_out0 = v_EQ_2591_out0;
assign v_EQ_3822_out0 = v_EQ_2592_out0;
assign v__10652_out0 = { v__4550_out0,v_S_8905_out0 };
assign v__10667_out0 = { v__4565_out0,v_S_9369_out0 };
assign v_MI_10833_out0 = v_MI_560_out0;
assign v_MI_10834_out0 = v_MI_561_out0;
assign v_JMIN_2662_out0 = v_MI_10833_out0;
assign v_JMIN_2663_out0 = v_MI_10834_out0;
assign v_JEQZ_10514_out0 = v_EQ_3821_out0;
assign v_JEQZ_10515_out0 = v_EQ_3822_out0;
assign v__10947_out0 = { v__10652_out0,v_CARRY_4904_out0 };
assign v__10962_out0 = { v__10667_out0,v_CARRY_5368_out0 };
assign v_JMIN_1205_out0 = v_JMIN_2662_out0;
assign v_JMIN_1206_out0 = v_JMIN_2663_out0;
assign v_JEQZ_2981_out0 = v_JEQZ_10514_out0;
assign v_JEQZ_2982_out0 = v_JEQZ_10515_out0;
assign v_COUT_10917_out0 = v__10947_out0;
assign v_COUT_10932_out0 = v__10962_out0;
assign v_CIN_2357_out0 = v_COUT_10917_out0;
assign v_CIN_2372_out0 = v_COUT_10932_out0;
assign v_G4_4846_out0 = v_JEQZ_2981_out0 && v_JEQ_8806_out0;
assign v_G4_4847_out0 = v_JEQZ_2982_out0 && v_JEQ_8807_out0;
assign v_G5_10533_out0 = v_JMIN_1205_out0 && v_JMI_3212_out0;
assign v_G5_10534_out0 = v_JMIN_1206_out0 && v_JMI_3213_out0;
assign v__470_out0 = v_CIN_2357_out0[8:8];
assign v__485_out0 = v_CIN_2372_out0[8:8];
assign v__1775_out0 = v_CIN_2357_out0[6:6];
assign v__1790_out0 = v_CIN_2372_out0[6:6];
assign v__2157_out0 = v_CIN_2357_out0[3:3];
assign v__2172_out0 = v_CIN_2372_out0[3:3];
assign v__2196_out0 = v_CIN_2357_out0[15:15];
assign v__2210_out0 = v_CIN_2372_out0[15:15];
assign v__2504_out0 = v_CIN_2357_out0[0:0];
assign v__2519_out0 = v_CIN_2372_out0[0:0];
assign v__3053_out0 = v_CIN_2357_out0[9:9];
assign v__3068_out0 = v_CIN_2372_out0[9:9];
assign v__3087_out0 = v_CIN_2357_out0[2:2];
assign v__3102_out0 = v_CIN_2372_out0[2:2];
assign v__3141_out0 = v_CIN_2357_out0[7:7];
assign v__3156_out0 = v_CIN_2372_out0[7:7];
assign v__3825_out0 = v_CIN_2357_out0[1:1];
assign v__3840_out0 = v_CIN_2372_out0[1:1];
assign v__3863_out0 = v_CIN_2357_out0[10:10];
assign v__3878_out0 = v_CIN_2372_out0[10:10];
assign v__6802_out0 = v_CIN_2357_out0[11:11];
assign v__6817_out0 = v_CIN_2372_out0[11:11];
assign v__7646_out0 = v_CIN_2357_out0[12:12];
assign v__7661_out0 = v_CIN_2372_out0[12:12];
assign v__8701_out0 = v_CIN_2357_out0[13:13];
assign v__8716_out0 = v_CIN_2372_out0[13:13];
assign v__8771_out0 = v_CIN_2357_out0[14:14];
assign v__8786_out0 = v_CIN_2372_out0[14:14];
assign v__10721_out0 = v_CIN_2357_out0[5:5];
assign v__10736_out0 = v_CIN_2372_out0[5:5];
assign v__13450_out0 = v_CIN_2357_out0[4:4];
assign v__13465_out0 = v_CIN_2372_out0[4:4];
assign v_G2_13645_out0 = v_JMP_546_out0 || v_G5_10533_out0;
assign v_G2_13646_out0 = v_JMP_547_out0 || v_G5_10534_out0;
assign v_RM_3384_out0 = v__7646_out0;
assign v_RM_3385_out0 = v__8771_out0;
assign v_RM_3387_out0 = v__10721_out0;
assign v_RM_3388_out0 = v__13450_out0;
assign v_RM_3389_out0 = v__8701_out0;
assign v_RM_3390_out0 = v__3053_out0;
assign v_RM_3391_out0 = v__3863_out0;
assign v_RM_3392_out0 = v__3825_out0;
assign v_RM_3393_out0 = v__2157_out0;
assign v_RM_3394_out0 = v__1775_out0;
assign v_RM_3395_out0 = v__3141_out0;
assign v_RM_3396_out0 = v__6802_out0;
assign v_RM_3397_out0 = v__470_out0;
assign v_RM_3398_out0 = v__3087_out0;
assign v_RM_3608_out0 = v__7661_out0;
assign v_RM_3609_out0 = v__8786_out0;
assign v_RM_3611_out0 = v__10736_out0;
assign v_RM_3612_out0 = v__13465_out0;
assign v_RM_3613_out0 = v__8716_out0;
assign v_RM_3614_out0 = v__3068_out0;
assign v_RM_3615_out0 = v__3878_out0;
assign v_RM_3616_out0 = v__3840_out0;
assign v_RM_3617_out0 = v__2172_out0;
assign v_RM_3618_out0 = v__1790_out0;
assign v_RM_3619_out0 = v__3156_out0;
assign v_RM_3620_out0 = v__6817_out0;
assign v_RM_3621_out0 = v__485_out0;
assign v_RM_3622_out0 = v__3102_out0;
assign v_G3_3812_out0 = v_G2_13645_out0 || v_G4_4846_out0;
assign v_G3_3813_out0 = v_G2_13646_out0 || v_G4_4847_out0;
assign v_CIN_9839_out0 = v__2196_out0;
assign v_CIN_10063_out0 = v__2210_out0;
assign v_RM_11375_out0 = v__2504_out0;
assign v_RM_11839_out0 = v__2519_out0;
assign v_JUMP_2187_out0 = v_G3_3812_out0;
assign v_JUMP_2188_out0 = v_G3_3813_out0;
assign v_RD_5928_out0 = v_CIN_9839_out0;
assign v_RD_6392_out0 = v_CIN_10063_out0;
assign v_G1_7790_out0 = ((v_RD_5935_out0 && !v_RM_11375_out0) || (!v_RD_5935_out0) && v_RM_11375_out0);
assign v_G1_8254_out0 = ((v_RD_6399_out0 && !v_RM_11839_out0) || (!v_RD_6399_out0) && v_RM_11839_out0);
assign v_RM_11363_out0 = v_RM_3384_out0;
assign v_RM_11365_out0 = v_RM_3385_out0;
assign v_RM_11369_out0 = v_RM_3387_out0;
assign v_RM_11371_out0 = v_RM_3388_out0;
assign v_RM_11373_out0 = v_RM_3389_out0;
assign v_RM_11376_out0 = v_RM_3390_out0;
assign v_RM_11378_out0 = v_RM_3391_out0;
assign v_RM_11380_out0 = v_RM_3392_out0;
assign v_RM_11382_out0 = v_RM_3393_out0;
assign v_RM_11384_out0 = v_RM_3394_out0;
assign v_RM_11386_out0 = v_RM_3395_out0;
assign v_RM_11388_out0 = v_RM_3396_out0;
assign v_RM_11390_out0 = v_RM_3397_out0;
assign v_RM_11392_out0 = v_RM_3398_out0;
assign v_RM_11827_out0 = v_RM_3608_out0;
assign v_RM_11829_out0 = v_RM_3609_out0;
assign v_RM_11833_out0 = v_RM_3611_out0;
assign v_RM_11835_out0 = v_RM_3612_out0;
assign v_RM_11837_out0 = v_RM_3613_out0;
assign v_RM_11840_out0 = v_RM_3614_out0;
assign v_RM_11842_out0 = v_RM_3615_out0;
assign v_RM_11844_out0 = v_RM_3616_out0;
assign v_RM_11846_out0 = v_RM_3617_out0;
assign v_RM_11848_out0 = v_RM_3618_out0;
assign v_RM_11850_out0 = v_RM_3619_out0;
assign v_RM_11852_out0 = v_RM_3620_out0;
assign v_RM_11854_out0 = v_RM_3621_out0;
assign v_RM_11856_out0 = v_RM_3622_out0;
assign v_G2_12326_out0 = v_RD_5935_out0 && v_RM_11375_out0;
assign v_G2_12790_out0 = v_RD_6399_out0 && v_RM_11839_out0;
assign v_G14_1178_out0 = v_G15_1855_out0 && v_JUMP_2187_out0;
assign v_G14_1179_out0 = v_G15_1856_out0 && v_JUMP_2188_out0;
assign v_CARRY_4935_out0 = v_G2_12326_out0;
assign v_CARRY_5399_out0 = v_G2_12790_out0;
assign v_G1_7778_out0 = ((v_RD_5923_out0 && !v_RM_11363_out0) || (!v_RD_5923_out0) && v_RM_11363_out0);
assign v_G1_7780_out0 = ((v_RD_5925_out0 && !v_RM_11365_out0) || (!v_RD_5925_out0) && v_RM_11365_out0);
assign v_G1_7784_out0 = ((v_RD_5929_out0 && !v_RM_11369_out0) || (!v_RD_5929_out0) && v_RM_11369_out0);
assign v_G1_7786_out0 = ((v_RD_5931_out0 && !v_RM_11371_out0) || (!v_RD_5931_out0) && v_RM_11371_out0);
assign v_G1_7788_out0 = ((v_RD_5933_out0 && !v_RM_11373_out0) || (!v_RD_5933_out0) && v_RM_11373_out0);
assign v_G1_7791_out0 = ((v_RD_5936_out0 && !v_RM_11376_out0) || (!v_RD_5936_out0) && v_RM_11376_out0);
assign v_G1_7793_out0 = ((v_RD_5938_out0 && !v_RM_11378_out0) || (!v_RD_5938_out0) && v_RM_11378_out0);
assign v_G1_7795_out0 = ((v_RD_5940_out0 && !v_RM_11380_out0) || (!v_RD_5940_out0) && v_RM_11380_out0);
assign v_G1_7797_out0 = ((v_RD_5942_out0 && !v_RM_11382_out0) || (!v_RD_5942_out0) && v_RM_11382_out0);
assign v_G1_7799_out0 = ((v_RD_5944_out0 && !v_RM_11384_out0) || (!v_RD_5944_out0) && v_RM_11384_out0);
assign v_G1_7801_out0 = ((v_RD_5946_out0 && !v_RM_11386_out0) || (!v_RD_5946_out0) && v_RM_11386_out0);
assign v_G1_7803_out0 = ((v_RD_5948_out0 && !v_RM_11388_out0) || (!v_RD_5948_out0) && v_RM_11388_out0);
assign v_G1_7805_out0 = ((v_RD_5950_out0 && !v_RM_11390_out0) || (!v_RD_5950_out0) && v_RM_11390_out0);
assign v_G1_7807_out0 = ((v_RD_5952_out0 && !v_RM_11392_out0) || (!v_RD_5952_out0) && v_RM_11392_out0);
assign v_G1_8242_out0 = ((v_RD_6387_out0 && !v_RM_11827_out0) || (!v_RD_6387_out0) && v_RM_11827_out0);
assign v_G1_8244_out0 = ((v_RD_6389_out0 && !v_RM_11829_out0) || (!v_RD_6389_out0) && v_RM_11829_out0);
assign v_G1_8248_out0 = ((v_RD_6393_out0 && !v_RM_11833_out0) || (!v_RD_6393_out0) && v_RM_11833_out0);
assign v_G1_8250_out0 = ((v_RD_6395_out0 && !v_RM_11835_out0) || (!v_RD_6395_out0) && v_RM_11835_out0);
assign v_G1_8252_out0 = ((v_RD_6397_out0 && !v_RM_11837_out0) || (!v_RD_6397_out0) && v_RM_11837_out0);
assign v_G1_8255_out0 = ((v_RD_6400_out0 && !v_RM_11840_out0) || (!v_RD_6400_out0) && v_RM_11840_out0);
assign v_G1_8257_out0 = ((v_RD_6402_out0 && !v_RM_11842_out0) || (!v_RD_6402_out0) && v_RM_11842_out0);
assign v_G1_8259_out0 = ((v_RD_6404_out0 && !v_RM_11844_out0) || (!v_RD_6404_out0) && v_RM_11844_out0);
assign v_G1_8261_out0 = ((v_RD_6406_out0 && !v_RM_11846_out0) || (!v_RD_6406_out0) && v_RM_11846_out0);
assign v_G1_8263_out0 = ((v_RD_6408_out0 && !v_RM_11848_out0) || (!v_RD_6408_out0) && v_RM_11848_out0);
assign v_G1_8265_out0 = ((v_RD_6410_out0 && !v_RM_11850_out0) || (!v_RD_6410_out0) && v_RM_11850_out0);
assign v_G1_8267_out0 = ((v_RD_6412_out0 && !v_RM_11852_out0) || (!v_RD_6412_out0) && v_RM_11852_out0);
assign v_G1_8269_out0 = ((v_RD_6414_out0 && !v_RM_11854_out0) || (!v_RD_6414_out0) && v_RM_11854_out0);
assign v_G1_8271_out0 = ((v_RD_6416_out0 && !v_RM_11856_out0) || (!v_RD_6416_out0) && v_RM_11856_out0);
assign v_S_8936_out0 = v_G1_7790_out0;
assign v_S_9400_out0 = v_G1_8254_out0;
assign v_G2_12314_out0 = v_RD_5923_out0 && v_RM_11363_out0;
assign v_G2_12316_out0 = v_RD_5925_out0 && v_RM_11365_out0;
assign v_G2_12320_out0 = v_RD_5929_out0 && v_RM_11369_out0;
assign v_G2_12322_out0 = v_RD_5931_out0 && v_RM_11371_out0;
assign v_G2_12324_out0 = v_RD_5933_out0 && v_RM_11373_out0;
assign v_G2_12327_out0 = v_RD_5936_out0 && v_RM_11376_out0;
assign v_G2_12329_out0 = v_RD_5938_out0 && v_RM_11378_out0;
assign v_G2_12331_out0 = v_RD_5940_out0 && v_RM_11380_out0;
assign v_G2_12333_out0 = v_RD_5942_out0 && v_RM_11382_out0;
assign v_G2_12335_out0 = v_RD_5944_out0 && v_RM_11384_out0;
assign v_G2_12337_out0 = v_RD_5946_out0 && v_RM_11386_out0;
assign v_G2_12339_out0 = v_RD_5948_out0 && v_RM_11388_out0;
assign v_G2_12341_out0 = v_RD_5950_out0 && v_RM_11390_out0;
assign v_G2_12343_out0 = v_RD_5952_out0 && v_RM_11392_out0;
assign v_G2_12778_out0 = v_RD_6387_out0 && v_RM_11827_out0;
assign v_G2_12780_out0 = v_RD_6389_out0 && v_RM_11829_out0;
assign v_G2_12784_out0 = v_RD_6393_out0 && v_RM_11833_out0;
assign v_G2_12786_out0 = v_RD_6395_out0 && v_RM_11835_out0;
assign v_G2_12788_out0 = v_RD_6397_out0 && v_RM_11837_out0;
assign v_G2_12791_out0 = v_RD_6400_out0 && v_RM_11840_out0;
assign v_G2_12793_out0 = v_RD_6402_out0 && v_RM_11842_out0;
assign v_G2_12795_out0 = v_RD_6404_out0 && v_RM_11844_out0;
assign v_G2_12797_out0 = v_RD_6406_out0 && v_RM_11846_out0;
assign v_G2_12799_out0 = v_RD_6408_out0 && v_RM_11848_out0;
assign v_G2_12801_out0 = v_RD_6410_out0 && v_RM_11850_out0;
assign v_G2_12803_out0 = v_RD_6412_out0 && v_RM_11852_out0;
assign v_G2_12805_out0 = v_RD_6414_out0 && v_RM_11854_out0;
assign v_G2_12807_out0 = v_RD_6416_out0 && v_RM_11856_out0;
assign v_S_4667_out0 = v_S_8936_out0;
assign v_S_4682_out0 = v_S_9400_out0;
assign v_CARRY_4923_out0 = v_G2_12314_out0;
assign v_CARRY_4925_out0 = v_G2_12316_out0;
assign v_CARRY_4929_out0 = v_G2_12320_out0;
assign v_CARRY_4931_out0 = v_G2_12322_out0;
assign v_CARRY_4933_out0 = v_G2_12324_out0;
assign v_CARRY_4936_out0 = v_G2_12327_out0;
assign v_CARRY_4938_out0 = v_G2_12329_out0;
assign v_CARRY_4940_out0 = v_G2_12331_out0;
assign v_CARRY_4942_out0 = v_G2_12333_out0;
assign v_CARRY_4944_out0 = v_G2_12335_out0;
assign v_CARRY_4946_out0 = v_G2_12337_out0;
assign v_CARRY_4948_out0 = v_G2_12339_out0;
assign v_CARRY_4950_out0 = v_G2_12341_out0;
assign v_CARRY_4952_out0 = v_G2_12343_out0;
assign v_CARRY_5387_out0 = v_G2_12778_out0;
assign v_CARRY_5389_out0 = v_G2_12780_out0;
assign v_CARRY_5393_out0 = v_G2_12784_out0;
assign v_CARRY_5395_out0 = v_G2_12786_out0;
assign v_CARRY_5397_out0 = v_G2_12788_out0;
assign v_CARRY_5400_out0 = v_G2_12791_out0;
assign v_CARRY_5402_out0 = v_G2_12793_out0;
assign v_CARRY_5404_out0 = v_G2_12795_out0;
assign v_CARRY_5406_out0 = v_G2_12797_out0;
assign v_CARRY_5408_out0 = v_G2_12799_out0;
assign v_CARRY_5410_out0 = v_G2_12801_out0;
assign v_CARRY_5412_out0 = v_G2_12803_out0;
assign v_CARRY_5414_out0 = v_G2_12805_out0;
assign v_CARRY_5416_out0 = v_G2_12807_out0;
assign v_S_8924_out0 = v_G1_7778_out0;
assign v_S_8926_out0 = v_G1_7780_out0;
assign v_S_8930_out0 = v_G1_7784_out0;
assign v_S_8932_out0 = v_G1_7786_out0;
assign v_S_8934_out0 = v_G1_7788_out0;
assign v_S_8937_out0 = v_G1_7791_out0;
assign v_S_8939_out0 = v_G1_7793_out0;
assign v_S_8941_out0 = v_G1_7795_out0;
assign v_S_8943_out0 = v_G1_7797_out0;
assign v_S_8945_out0 = v_G1_7799_out0;
assign v_S_8947_out0 = v_G1_7801_out0;
assign v_S_8949_out0 = v_G1_7803_out0;
assign v_S_8951_out0 = v_G1_7805_out0;
assign v_S_8953_out0 = v_G1_7807_out0;
assign v_S_9388_out0 = v_G1_8242_out0;
assign v_S_9390_out0 = v_G1_8244_out0;
assign v_S_9394_out0 = v_G1_8248_out0;
assign v_S_9396_out0 = v_G1_8250_out0;
assign v_S_9398_out0 = v_G1_8252_out0;
assign v_S_9401_out0 = v_G1_8255_out0;
assign v_S_9403_out0 = v_G1_8257_out0;
assign v_S_9405_out0 = v_G1_8259_out0;
assign v_S_9407_out0 = v_G1_8261_out0;
assign v_S_9409_out0 = v_G1_8263_out0;
assign v_S_9411_out0 = v_G1_8265_out0;
assign v_S_9413_out0 = v_G1_8267_out0;
assign v_S_9415_out0 = v_G1_8269_out0;
assign v_S_9417_out0 = v_G1_8271_out0;
assign v_CIN_9845_out0 = v_CARRY_4935_out0;
assign v_CIN_10069_out0 = v_CARRY_5399_out0;
assign v_MUX1_10773_out0 = v_G14_1178_out0 ? v_JUMPADRESS_4745_out0 : v_REG1_432_out0;
assign v_MUX1_10774_out0 = v_G14_1179_out0 ? v_JUMPADRESS_4746_out0 : v_REG1_433_out0;
assign v__1716_out0 = { v__3223_out0,v_S_4667_out0 };
assign v__1717_out0 = { v__3224_out0,v_S_4682_out0 };
assign v_RD_5941_out0 = v_CIN_9845_out0;
assign v_RD_6405_out0 = v_CIN_10069_out0;
assign {v_A1_7019_out1,v_A1_7019_out0 } = v_MUX1_10773_out0 + v_ADDER_IN_10995_out0 + v_G22_1899_out0;
assign {v_A1_7020_out1,v_A1_7020_out0 } = v_MUX1_10774_out0 + v_ADDER_IN_10996_out0 + v_G22_1900_out0;
assign v_RM_11364_out0 = v_S_8924_out0;
assign v_RM_11366_out0 = v_S_8926_out0;
assign v_RM_11370_out0 = v_S_8930_out0;
assign v_RM_11372_out0 = v_S_8932_out0;
assign v_RM_11374_out0 = v_S_8934_out0;
assign v_RM_11377_out0 = v_S_8937_out0;
assign v_RM_11379_out0 = v_S_8939_out0;
assign v_RM_11381_out0 = v_S_8941_out0;
assign v_RM_11383_out0 = v_S_8943_out0;
assign v_RM_11385_out0 = v_S_8945_out0;
assign v_RM_11387_out0 = v_S_8947_out0;
assign v_RM_11389_out0 = v_S_8949_out0;
assign v_RM_11391_out0 = v_S_8951_out0;
assign v_RM_11393_out0 = v_S_8953_out0;
assign v_RM_11828_out0 = v_S_9388_out0;
assign v_RM_11830_out0 = v_S_9390_out0;
assign v_RM_11834_out0 = v_S_9394_out0;
assign v_RM_11836_out0 = v_S_9396_out0;
assign v_RM_11838_out0 = v_S_9398_out0;
assign v_RM_11841_out0 = v_S_9401_out0;
assign v_RM_11843_out0 = v_S_9403_out0;
assign v_RM_11845_out0 = v_S_9405_out0;
assign v_RM_11847_out0 = v_S_9407_out0;
assign v_RM_11849_out0 = v_S_9409_out0;
assign v_RM_11851_out0 = v_S_9411_out0;
assign v_RM_11853_out0 = v_S_9413_out0;
assign v_RM_11855_out0 = v_S_9415_out0;
assign v_RM_11857_out0 = v_S_9417_out0;
assign v_COUT_70_out0 = v_A1_7019_out1;
assign v_COUT_71_out0 = v_A1_7020_out1;
assign v_G1_7796_out0 = ((v_RD_5941_out0 && !v_RM_11381_out0) || (!v_RD_5941_out0) && v_RM_11381_out0);
assign v_G1_8260_out0 = ((v_RD_6405_out0 && !v_RM_11845_out0) || (!v_RD_6405_out0) && v_RM_11845_out0);
assign v_MUX3_10330_out0 = v_STP_11240_out0 ? v_A1_7019_out0 : v_MUX1_10773_out0;
assign v_MUX3_10331_out0 = v_STP_11241_out0 ? v_A1_7020_out0 : v_MUX1_10774_out0;
assign v_MUX5_10845_out0 = v_STORE_WEN_4544_out0 ? v_REG1_432_out0 : v_A1_7019_out0;
assign v_MUX5_10846_out0 = v_STORE_WEN_4545_out0 ? v_REG1_433_out0 : v_A1_7020_out0;
assign v_G2_12332_out0 = v_RD_5941_out0 && v_RM_11381_out0;
assign v_G2_12796_out0 = v_RD_6405_out0 && v_RM_11845_out0;
assign v_MUX4_2658_out0 = v_BYTE_READY_2852_out0 ? v_C1_2426_out0 : v_MUX5_10845_out0;
assign v_MUX4_2659_out0 = v_BYTE_READY_2853_out0 ? v_C1_2427_out0 : v_MUX5_10846_out0;
assign v_CARRY_4941_out0 = v_G2_12332_out0;
assign v_CARRY_5405_out0 = v_G2_12796_out0;
assign v_PC_COUNTER_NEXT_7064_out0 = v_MUX3_10330_out0;
assign v_PC_COUNTER_NEXT_7065_out0 = v_MUX3_10331_out0;
assign v_S_8942_out0 = v_G1_7796_out0;
assign v_S_9406_out0 = v_G1_8260_out0;
assign v_PC_COUNTER_25_out0 = v_PC_COUNTER_NEXT_7064_out0;
assign v_PC_COUNTER_26_out0 = v_PC_COUNTER_NEXT_7065_out0;
assign v_REGISTER_216_out0 = v_MUX4_2658_out0;
assign v_REGISTER_217_out0 = v_MUX4_2659_out0;
assign v_S_1256_out0 = v_S_8942_out0;
assign v_S_1480_out0 = v_S_9406_out0;
assign v_G1_4032_out0 = v_CARRY_4941_out0 || v_CARRY_4940_out0;
assign v_G1_4256_out0 = v_CARRY_5405_out0 || v_CARRY_5404_out0;
assign v_COUT_724_out0 = v_G1_4032_out0;
assign v_COUT_948_out0 = v_G1_4256_out0;
assign v_MUX3_3225_out0 = v_BYTE_READY_7021_out0 ? v_C2_10761_out0 : v_PC_COUNTER_25_out0;
assign v_MUX3_3226_out0 = v_BYTE_READY_7022_out0 ? v_C2_10762_out0 : v_PC_COUNTER_26_out0;
assign v__8697_out0 = { v_PC_COUNTER_25_out0,v_C1_2005_out0 };
assign v__8698_out0 = { v_PC_COUNTER_26_out0,v_C1_2006_out0 };
assign v_REGISTER_13346_out0 = v_REGISTER_216_out0;
assign v_REGISTER_13347_out0 = v_REGISTER_217_out0;
assign v_REGISTER4_1705_out0 = v_REGISTER_13346_out0;
assign v_REGISTER4_1706_out0 = v_REGISTER_13347_out0;
assign v_MUX2_3202_out0 = v_BYTE_READY_7021_out0 ? v__8697_out0 : v_RAM_IN_233_out0;
assign v_MUX2_3203_out0 = v_BYTE_READY_7022_out0 ? v__8698_out0 : v_RAM_IN_234_out0;
assign v_CIN_9851_out0 = v_COUT_724_out0;
assign v_CIN_10075_out0 = v_COUT_948_out0;
assign v_NEXTADD_10526_out0 = v_MUX3_3225_out0;
assign v_NEXTADD_10527_out0 = v_MUX3_3226_out0;
assign v_NEXTADRESS_1803_out0 = v_NEXTADD_10526_out0;
assign v_NEXTADRESS_1804_out0 = v_NEXTADD_10527_out0;
assign v_REGISTER14_3201_out0 = v_REGISTER4_1706_out0;
assign v_RD_5953_out0 = v_CIN_9851_out0;
assign v_RD_6417_out0 = v_CIN_10075_out0;
assign v_REGISTER15_8833_out0 = v_REGISTER4_1705_out0;
assign v_DATA_IN_10552_out0 = v_MUX2_3202_out0;
assign v_DATA_IN_10553_out0 = v_MUX2_3203_out0;
assign v_DATA_RAM_IN_558_out0 = v_DATA_IN_10552_out0;
assign v_DATA_RAM_IN_559_out0 = v_DATA_IN_10553_out0;
assign v_NEXT_ADRESS_3243_out0 = v_NEXTADRESS_1803_out0;
assign v_NEXT_ADRESS_3244_out0 = v_NEXTADRESS_1804_out0;
assign v_G1_7808_out0 = ((v_RD_5953_out0 && !v_RM_11393_out0) || (!v_RD_5953_out0) && v_RM_11393_out0);
assign v_G1_8272_out0 = ((v_RD_6417_out0 && !v_RM_11857_out0) || (!v_RD_6417_out0) && v_RM_11857_out0);
assign v_G2_12344_out0 = v_RD_5953_out0 && v_RM_11393_out0;
assign v_G2_12808_out0 = v_RD_6417_out0 && v_RM_11857_out0;
assign v_DATA_RAM_IN0_284_out0 = v_DATA_RAM_IN_559_out0;
assign v_DATA_RAM_IN1_4779_out0 = v_DATA_RAM_IN_558_out0;
assign v_CARRY_4953_out0 = v_G2_12344_out0;
assign v_CARRY_5417_out0 = v_G2_12808_out0;
assign v_S_8954_out0 = v_G1_7808_out0;
assign v_S_9418_out0 = v_G1_8272_out0;
assign v_ADRESS_ins1_10617_out0 = v_NEXT_ADRESS_3243_out0;
assign v_ADRESS_ins0_11169_out0 = v_NEXT_ADRESS_3244_out0;
assign v_DATA1_603_out0 = v_DATA_RAM_IN1_4779_out0;
assign v_S_1262_out0 = v_S_8954_out0;
assign v_S_1486_out0 = v_S_9418_out0;
assign v_G1_4038_out0 = v_CARRY_4953_out0 || v_CARRY_4952_out0;
assign v_G1_4262_out0 = v_CARRY_5417_out0 || v_CARRY_5416_out0;
assign v_DATA0_4737_out0 = v_DATA_RAM_IN0_284_out0;
assign v_COUT_730_out0 = v_G1_4038_out0;
assign v_COUT_954_out0 = v_G1_4262_out0;
assign v_DATA1_1974_out0 = v_DATA1_603_out0;
assign v__4784_out0 = { v_S_1256_out0,v_S_1262_out0 };
assign v__4799_out0 = { v_S_1480_out0,v_S_1486_out0 };
assign v_DATA0_13293_out0 = v_DATA0_4737_out0;
assign v_MUX4_1698_out0 = v_TX_inst0_608_out0 ? v_DATA0_13293_out0 : v_DATA1_1974_out0;
assign v_CIN_9846_out0 = v_COUT_730_out0;
assign v_CIN_10070_out0 = v_COUT_954_out0;
assign v_MUX3_10787_out0 = v_MUX_ENABLE_2349_out0 ? v_DATA0_13293_out0 : v_DATA1_1974_out0;
assign v_DATA_to_transmit_4546_out0 = v_MUX4_1698_out0;
assign v_RD_5943_out0 = v_CIN_9846_out0;
assign v_RD_6407_out0 = v_CIN_10070_out0;
assign v_DATA_10445_out0 = v_MUX3_10787_out0;
assign v_DATA_2469_out0 = v_DATA_10445_out0;
assign v_REGISTER_OUTPUT_3268_out0 = v_DATA_to_transmit_4546_out0;
assign v_G1_7798_out0 = ((v_RD_5943_out0 && !v_RM_11383_out0) || (!v_RD_5943_out0) && v_RM_11383_out0);
assign v_G1_8262_out0 = ((v_RD_6407_out0 && !v_RM_11847_out0) || (!v_RD_6407_out0) && v_RM_11847_out0);
assign v_G2_12334_out0 = v_RD_5943_out0 && v_RM_11383_out0;
assign v_G2_12798_out0 = v_RD_6407_out0 && v_RM_11847_out0;
assign v_REGISTER_OUTPUT2_2398_out0 = v_REGISTER_OUTPUT_3268_out0;
assign v_CARRY_4943_out0 = v_G2_12334_out0;
assign v_CARRY_5407_out0 = v_G2_12798_out0;
assign v_S_8944_out0 = v_G1_7798_out0;
assign v_S_9408_out0 = v_G1_8262_out0;
assign v_S_1257_out0 = v_S_8944_out0;
assign v_S_1481_out0 = v_S_9408_out0;
assign v_split_3196_out0 = v_REGISTER_OUTPUT2_2398_out0[7:0];
assign v_split_3196_out1 = v_REGISTER_OUTPUT2_2398_out0[15:8];
assign v_G1_4033_out0 = v_CARRY_4943_out0 || v_CARRY_4942_out0;
assign v_G1_4257_out0 = v_CARRY_5407_out0 || v_CARRY_5406_out0;
assign v_COUT_725_out0 = v_G1_4033_out0;
assign v_COUT_949_out0 = v_G1_4257_out0;
assign v__2554_out0 = { v__4784_out0,v_S_1257_out0 };
assign v__2569_out0 = { v__4799_out0,v_S_1481_out0 };
assign v_MUX1_13260_out0 = v_BYTE_COMP_1_8743_out0 ? v_split_3196_out1 : v_split_3196_out0;
assign v_TRANSMISSION_DATA2_7014_out0 = v_MUX1_13260_out0;
assign v_CIN_9841_out0 = v_COUT_725_out0;
assign v_CIN_10065_out0 = v_COUT_949_out0;
assign v_REGISTER_TRANSMIT_DATA_12241_out0 = v_MUX1_13260_out0;
assign v_TRANSMIT_DATA_76_out0 = v_REGISTER_TRANSMIT_DATA_12241_out0;
assign v_RD_5932_out0 = v_CIN_9841_out0;
assign v_RD_6396_out0 = v_CIN_10065_out0;
assign v_TRANSIMISSION_DATA_10818_out0 = v_TRANSMISSION_DATA2_7014_out0;
assign v_SEL1_240_out0 = v_TRANSMIT_DATA_76_out0[6:6];
assign v_SEL1_1164_out0 = v_TRANSMIT_DATA_76_out0[2:2];
assign v_SEL1_1204_out0 = v_TRANSMIT_DATA_76_out0[4:4];
assign v_SEL1_2319_out0 = v_TRANSMIT_DATA_76_out0[0:0];
assign v_SEL1_2428_out0 = v_TRANSMIT_DATA_76_out0[5:5];
assign v_SEL1_4858_out0 = v_TRANSMIT_DATA_76_out0[3:3];
assign v_G1_7787_out0 = ((v_RD_5932_out0 && !v_RM_11372_out0) || (!v_RD_5932_out0) && v_RM_11372_out0);
assign v_G1_8251_out0 = ((v_RD_6396_out0 && !v_RM_11836_out0) || (!v_RD_6396_out0) && v_RM_11836_out0);
assign v_SEL1_10304_out0 = v_TRANSMIT_DATA_76_out0[1:1];
assign v_G2_12323_out0 = v_RD_5932_out0 && v_RM_11372_out0;
assign v_G2_12787_out0 = v_RD_6396_out0 && v_RM_11836_out0;
assign v_SEL1_13445_out0 = v_TRANSMIT_DATA_76_out0[7:7];
assign v_MUX1_2625_out0 = v_transmit_INSTRUCTION_2674_out0 ? v_SEL1_240_out0 : v_FF1_1955_out0;
assign v_MUX4_3219_out0 = v_transmit_INSTRUCTION_2674_out0 ? v_SEL1_4858_out0 : v_FF4_463_out0;
assign v_MUX2_4448_out0 = v_transmit_INSTRUCTION_2674_out0 ? v_SEL1_2428_out0 : v_FF2_2833_out0;
assign v_CARRY_4932_out0 = v_G2_12323_out0;
assign v_CARRY_5396_out0 = v_G2_12787_out0;
assign v_MUX3_7140_out0 = v_transmit_INSTRUCTION_2674_out0 ? v_SEL1_1204_out0 : v_FF3_11046_out0;
assign v_S_8933_out0 = v_G1_7787_out0;
assign v_S_9397_out0 = v_G1_8251_out0;
assign v_MUX7_10448_out0 = v_transmit_INSTRUCTION_2674_out0 ? v_SEL1_2319_out0 : v_FF7_4781_out0;
assign v_MUX6_10976_out0 = v_transmit_INSTRUCTION_2674_out0 ? v_SEL1_10304_out0 : v_FF6_112_out0;
assign v_MUX5_13348_out0 = v_transmit_INSTRUCTION_2674_out0 ? v_SEL1_1164_out0 : v_FF5_7100_out0;
assign v_S_1252_out0 = v_S_8933_out0;
assign v_S_1476_out0 = v_S_9397_out0;
assign v_G1_4028_out0 = v_CARRY_4932_out0 || v_CARRY_4931_out0;
assign v_G1_4252_out0 = v_CARRY_5396_out0 || v_CARRY_5395_out0;
assign v_COUT_720_out0 = v_G1_4028_out0;
assign v_COUT_944_out0 = v_G1_4252_out0;
assign v__7034_out0 = { v__2554_out0,v_S_1252_out0 };
assign v__7049_out0 = { v__2569_out0,v_S_1476_out0 };
assign v_CIN_9840_out0 = v_COUT_720_out0;
assign v_CIN_10064_out0 = v_COUT_944_out0;
assign v_RD_5930_out0 = v_CIN_9840_out0;
assign v_RD_6394_out0 = v_CIN_10064_out0;
assign v_G1_7785_out0 = ((v_RD_5930_out0 && !v_RM_11370_out0) || (!v_RD_5930_out0) && v_RM_11370_out0);
assign v_G1_8249_out0 = ((v_RD_6394_out0 && !v_RM_11834_out0) || (!v_RD_6394_out0) && v_RM_11834_out0);
assign v_G2_12321_out0 = v_RD_5930_out0 && v_RM_11370_out0;
assign v_G2_12785_out0 = v_RD_6394_out0 && v_RM_11834_out0;
assign v_CARRY_4930_out0 = v_G2_12321_out0;
assign v_CARRY_5394_out0 = v_G2_12785_out0;
assign v_S_8931_out0 = v_G1_7785_out0;
assign v_S_9395_out0 = v_G1_8249_out0;
assign v_S_1251_out0 = v_S_8931_out0;
assign v_S_1475_out0 = v_S_9395_out0;
assign v_G1_4027_out0 = v_CARRY_4930_out0 || v_CARRY_4929_out0;
assign v_G1_4251_out0 = v_CARRY_5394_out0 || v_CARRY_5393_out0;
assign v_COUT_719_out0 = v_G1_4027_out0;
assign v_COUT_943_out0 = v_G1_4251_out0;
assign v__13520_out0 = { v__7034_out0,v_S_1251_out0 };
assign v__13535_out0 = { v__7049_out0,v_S_1475_out0 };
assign v_CIN_9847_out0 = v_COUT_719_out0;
assign v_CIN_10071_out0 = v_COUT_943_out0;
assign v_RD_5945_out0 = v_CIN_9847_out0;
assign v_RD_6409_out0 = v_CIN_10071_out0;
assign v_G1_7800_out0 = ((v_RD_5945_out0 && !v_RM_11385_out0) || (!v_RD_5945_out0) && v_RM_11385_out0);
assign v_G1_8264_out0 = ((v_RD_6409_out0 && !v_RM_11849_out0) || (!v_RD_6409_out0) && v_RM_11849_out0);
assign v_G2_12336_out0 = v_RD_5945_out0 && v_RM_11385_out0;
assign v_G2_12800_out0 = v_RD_6409_out0 && v_RM_11849_out0;
assign v_CARRY_4945_out0 = v_G2_12336_out0;
assign v_CARRY_5409_out0 = v_G2_12800_out0;
assign v_S_8946_out0 = v_G1_7800_out0;
assign v_S_9410_out0 = v_G1_8264_out0;
assign v_S_1258_out0 = v_S_8946_out0;
assign v_S_1482_out0 = v_S_9410_out0;
assign v_G1_4034_out0 = v_CARRY_4945_out0 || v_CARRY_4944_out0;
assign v_G1_4258_out0 = v_CARRY_5409_out0 || v_CARRY_5408_out0;
assign v_COUT_726_out0 = v_G1_4034_out0;
assign v_COUT_950_out0 = v_G1_4258_out0;
assign v__3313_out0 = { v__13520_out0,v_S_1258_out0 };
assign v__3328_out0 = { v__13535_out0,v_S_1482_out0 };
assign v_CIN_9848_out0 = v_COUT_726_out0;
assign v_CIN_10072_out0 = v_COUT_950_out0;
assign v_RD_5947_out0 = v_CIN_9848_out0;
assign v_RD_6411_out0 = v_CIN_10072_out0;
assign v_G1_7802_out0 = ((v_RD_5947_out0 && !v_RM_11387_out0) || (!v_RD_5947_out0) && v_RM_11387_out0);
assign v_G1_8266_out0 = ((v_RD_6411_out0 && !v_RM_11851_out0) || (!v_RD_6411_out0) && v_RM_11851_out0);
assign v_G2_12338_out0 = v_RD_5947_out0 && v_RM_11387_out0;
assign v_G2_12802_out0 = v_RD_6411_out0 && v_RM_11851_out0;
assign v_CARRY_4947_out0 = v_G2_12338_out0;
assign v_CARRY_5411_out0 = v_G2_12802_out0;
assign v_S_8948_out0 = v_G1_7802_out0;
assign v_S_9412_out0 = v_G1_8266_out0;
assign v_S_1259_out0 = v_S_8948_out0;
assign v_S_1483_out0 = v_S_9412_out0;
assign v_G1_4035_out0 = v_CARRY_4947_out0 || v_CARRY_4946_out0;
assign v_G1_4259_out0 = v_CARRY_5411_out0 || v_CARRY_5410_out0;
assign v_COUT_727_out0 = v_G1_4035_out0;
assign v_COUT_951_out0 = v_G1_4259_out0;
assign v__7149_out0 = { v__3313_out0,v_S_1259_out0 };
assign v__7164_out0 = { v__3328_out0,v_S_1483_out0 };
assign v_CIN_9850_out0 = v_COUT_727_out0;
assign v_CIN_10074_out0 = v_COUT_951_out0;
assign v_RD_5951_out0 = v_CIN_9850_out0;
assign v_RD_6415_out0 = v_CIN_10074_out0;
assign v_G1_7806_out0 = ((v_RD_5951_out0 && !v_RM_11391_out0) || (!v_RD_5951_out0) && v_RM_11391_out0);
assign v_G1_8270_out0 = ((v_RD_6415_out0 && !v_RM_11855_out0) || (!v_RD_6415_out0) && v_RM_11855_out0);
assign v_G2_12342_out0 = v_RD_5951_out0 && v_RM_11391_out0;
assign v_G2_12806_out0 = v_RD_6415_out0 && v_RM_11855_out0;
assign v_CARRY_4951_out0 = v_G2_12342_out0;
assign v_CARRY_5415_out0 = v_G2_12806_out0;
assign v_S_8952_out0 = v_G1_7806_out0;
assign v_S_9416_out0 = v_G1_8270_out0;
assign v_S_1261_out0 = v_S_8952_out0;
assign v_S_1485_out0 = v_S_9416_out0;
assign v_G1_4037_out0 = v_CARRY_4951_out0 || v_CARRY_4950_out0;
assign v_G1_4261_out0 = v_CARRY_5415_out0 || v_CARRY_5414_out0;
assign v_COUT_729_out0 = v_G1_4037_out0;
assign v_COUT_953_out0 = v_G1_4261_out0;
assign v__4751_out0 = { v__7149_out0,v_S_1261_out0 };
assign v__4766_out0 = { v__7164_out0,v_S_1485_out0 };
assign v_CIN_9843_out0 = v_COUT_729_out0;
assign v_CIN_10067_out0 = v_COUT_953_out0;
assign v_RD_5937_out0 = v_CIN_9843_out0;
assign v_RD_6401_out0 = v_CIN_10067_out0;
assign v_G1_7792_out0 = ((v_RD_5937_out0 && !v_RM_11377_out0) || (!v_RD_5937_out0) && v_RM_11377_out0);
assign v_G1_8256_out0 = ((v_RD_6401_out0 && !v_RM_11841_out0) || (!v_RD_6401_out0) && v_RM_11841_out0);
assign v_G2_12328_out0 = v_RD_5937_out0 && v_RM_11377_out0;
assign v_G2_12792_out0 = v_RD_6401_out0 && v_RM_11841_out0;
assign v_CARRY_4937_out0 = v_G2_12328_out0;
assign v_CARRY_5401_out0 = v_G2_12792_out0;
assign v_S_8938_out0 = v_G1_7792_out0;
assign v_S_9402_out0 = v_G1_8256_out0;
assign v_S_1254_out0 = v_S_8938_out0;
assign v_S_1478_out0 = v_S_9402_out0;
assign v_G1_4030_out0 = v_CARRY_4937_out0 || v_CARRY_4936_out0;
assign v_G1_4254_out0 = v_CARRY_5401_out0 || v_CARRY_5400_out0;
assign v_COUT_722_out0 = v_G1_4030_out0;
assign v_COUT_946_out0 = v_G1_4254_out0;
assign v__6928_out0 = { v__4751_out0,v_S_1254_out0 };
assign v__6943_out0 = { v__4766_out0,v_S_1478_out0 };
assign v_CIN_9844_out0 = v_COUT_722_out0;
assign v_CIN_10068_out0 = v_COUT_946_out0;
assign v_RD_5939_out0 = v_CIN_9844_out0;
assign v_RD_6403_out0 = v_CIN_10068_out0;
assign v_G1_7794_out0 = ((v_RD_5939_out0 && !v_RM_11379_out0) || (!v_RD_5939_out0) && v_RM_11379_out0);
assign v_G1_8258_out0 = ((v_RD_6403_out0 && !v_RM_11843_out0) || (!v_RD_6403_out0) && v_RM_11843_out0);
assign v_G2_12330_out0 = v_RD_5939_out0 && v_RM_11379_out0;
assign v_G2_12794_out0 = v_RD_6403_out0 && v_RM_11843_out0;
assign v_CARRY_4939_out0 = v_G2_12330_out0;
assign v_CARRY_5403_out0 = v_G2_12794_out0;
assign v_S_8940_out0 = v_G1_7794_out0;
assign v_S_9404_out0 = v_G1_8258_out0;
assign v_S_1255_out0 = v_S_8940_out0;
assign v_S_1479_out0 = v_S_9404_out0;
assign v_G1_4031_out0 = v_CARRY_4939_out0 || v_CARRY_4938_out0;
assign v_G1_4255_out0 = v_CARRY_5403_out0 || v_CARRY_5402_out0;
assign v_COUT_723_out0 = v_G1_4031_out0;
assign v_COUT_947_out0 = v_G1_4255_out0;
assign v__5804_out0 = { v__6928_out0,v_S_1255_out0 };
assign v__5819_out0 = { v__6943_out0,v_S_1479_out0 };
assign v_CIN_9849_out0 = v_COUT_723_out0;
assign v_CIN_10073_out0 = v_COUT_947_out0;
assign v_RD_5949_out0 = v_CIN_9849_out0;
assign v_RD_6413_out0 = v_CIN_10073_out0;
assign v_G1_7804_out0 = ((v_RD_5949_out0 && !v_RM_11389_out0) || (!v_RD_5949_out0) && v_RM_11389_out0);
assign v_G1_8268_out0 = ((v_RD_6413_out0 && !v_RM_11853_out0) || (!v_RD_6413_out0) && v_RM_11853_out0);
assign v_G2_12340_out0 = v_RD_5949_out0 && v_RM_11389_out0;
assign v_G2_12804_out0 = v_RD_6413_out0 && v_RM_11853_out0;
assign v_CARRY_4949_out0 = v_G2_12340_out0;
assign v_CARRY_5413_out0 = v_G2_12804_out0;
assign v_S_8950_out0 = v_G1_7804_out0;
assign v_S_9414_out0 = v_G1_8268_out0;
assign v_S_1260_out0 = v_S_8950_out0;
assign v_S_1484_out0 = v_S_9414_out0;
assign v_G1_4036_out0 = v_CARRY_4949_out0 || v_CARRY_4948_out0;
assign v_G1_4260_out0 = v_CARRY_5413_out0 || v_CARRY_5412_out0;
assign v_COUT_728_out0 = v_G1_4036_out0;
assign v_COUT_952_out0 = v_G1_4260_out0;
assign v__2028_out0 = { v__5804_out0,v_S_1260_out0 };
assign v__2043_out0 = { v__5819_out0,v_S_1484_out0 };
assign v_CIN_9837_out0 = v_COUT_728_out0;
assign v_CIN_10061_out0 = v_COUT_952_out0;
assign v_RD_5924_out0 = v_CIN_9837_out0;
assign v_RD_6388_out0 = v_CIN_10061_out0;
assign v_G1_7779_out0 = ((v_RD_5924_out0 && !v_RM_11364_out0) || (!v_RD_5924_out0) && v_RM_11364_out0);
assign v_G1_8243_out0 = ((v_RD_6388_out0 && !v_RM_11828_out0) || (!v_RD_6388_out0) && v_RM_11828_out0);
assign v_G2_12315_out0 = v_RD_5924_out0 && v_RM_11364_out0;
assign v_G2_12779_out0 = v_RD_6388_out0 && v_RM_11828_out0;
assign v_CARRY_4924_out0 = v_G2_12315_out0;
assign v_CARRY_5388_out0 = v_G2_12779_out0;
assign v_S_8925_out0 = v_G1_7779_out0;
assign v_S_9389_out0 = v_G1_8243_out0;
assign v_S_1248_out0 = v_S_8925_out0;
assign v_S_1472_out0 = v_S_9389_out0;
assign v_G1_4024_out0 = v_CARRY_4924_out0 || v_CARRY_4923_out0;
assign v_G1_4248_out0 = v_CARRY_5388_out0 || v_CARRY_5387_out0;
assign v_COUT_716_out0 = v_G1_4024_out0;
assign v_COUT_940_out0 = v_G1_4248_out0;
assign v__2795_out0 = { v__2028_out0,v_S_1248_out0 };
assign v__2810_out0 = { v__2043_out0,v_S_1472_out0 };
assign v_CIN_9842_out0 = v_COUT_716_out0;
assign v_CIN_10066_out0 = v_COUT_940_out0;
assign v_RD_5934_out0 = v_CIN_9842_out0;
assign v_RD_6398_out0 = v_CIN_10066_out0;
assign v_G1_7789_out0 = ((v_RD_5934_out0 && !v_RM_11374_out0) || (!v_RD_5934_out0) && v_RM_11374_out0);
assign v_G1_8253_out0 = ((v_RD_6398_out0 && !v_RM_11838_out0) || (!v_RD_6398_out0) && v_RM_11838_out0);
assign v_G2_12325_out0 = v_RD_5934_out0 && v_RM_11374_out0;
assign v_G2_12789_out0 = v_RD_6398_out0 && v_RM_11838_out0;
assign v_CARRY_4934_out0 = v_G2_12325_out0;
assign v_CARRY_5398_out0 = v_G2_12789_out0;
assign v_S_8935_out0 = v_G1_7789_out0;
assign v_S_9399_out0 = v_G1_8253_out0;
assign v_S_1253_out0 = v_S_8935_out0;
assign v_S_1477_out0 = v_S_9399_out0;
assign v_G1_4029_out0 = v_CARRY_4934_out0 || v_CARRY_4933_out0;
assign v_G1_4253_out0 = v_CARRY_5398_out0 || v_CARRY_5397_out0;
assign v_COUT_721_out0 = v_G1_4029_out0;
assign v_COUT_945_out0 = v_G1_4253_out0;
assign v__1827_out0 = { v__2795_out0,v_S_1253_out0 };
assign v__1842_out0 = { v__2810_out0,v_S_1477_out0 };
assign v_CIN_9838_out0 = v_COUT_721_out0;
assign v_CIN_10062_out0 = v_COUT_945_out0;
assign v_RD_5926_out0 = v_CIN_9838_out0;
assign v_RD_6390_out0 = v_CIN_10062_out0;
assign v_G1_7781_out0 = ((v_RD_5926_out0 && !v_RM_11366_out0) || (!v_RD_5926_out0) && v_RM_11366_out0);
assign v_G1_8245_out0 = ((v_RD_6390_out0 && !v_RM_11830_out0) || (!v_RD_6390_out0) && v_RM_11830_out0);
assign v_G2_12317_out0 = v_RD_5926_out0 && v_RM_11366_out0;
assign v_G2_12781_out0 = v_RD_6390_out0 && v_RM_11830_out0;
assign v_CARRY_4926_out0 = v_G2_12317_out0;
assign v_CARRY_5390_out0 = v_G2_12781_out0;
assign v_S_8927_out0 = v_G1_7781_out0;
assign v_S_9391_out0 = v_G1_8245_out0;
assign v_S_1249_out0 = v_S_8927_out0;
assign v_S_1473_out0 = v_S_9391_out0;
assign v_G1_4025_out0 = v_CARRY_4926_out0 || v_CARRY_4925_out0;
assign v_G1_4249_out0 = v_CARRY_5390_out0 || v_CARRY_5389_out0;
assign v_COUT_717_out0 = v_G1_4025_out0;
assign v_COUT_941_out0 = v_G1_4249_out0;
assign v__4551_out0 = { v__1827_out0,v_S_1249_out0 };
assign v__4566_out0 = { v__1842_out0,v_S_1473_out0 };
assign v_RM_3386_out0 = v_COUT_717_out0;
assign v_RM_3610_out0 = v_COUT_941_out0;
assign v_RM_11367_out0 = v_RM_3386_out0;
assign v_RM_11831_out0 = v_RM_3610_out0;
assign v_G1_7782_out0 = ((v_RD_5927_out0 && !v_RM_11367_out0) || (!v_RD_5927_out0) && v_RM_11367_out0);
assign v_G1_8246_out0 = ((v_RD_6391_out0 && !v_RM_11831_out0) || (!v_RD_6391_out0) && v_RM_11831_out0);
assign v_G2_12318_out0 = v_RD_5927_out0 && v_RM_11367_out0;
assign v_G2_12782_out0 = v_RD_6391_out0 && v_RM_11831_out0;
assign v_CARRY_4927_out0 = v_G2_12318_out0;
assign v_CARRY_5391_out0 = v_G2_12782_out0;
assign v_S_8928_out0 = v_G1_7782_out0;
assign v_S_9392_out0 = v_G1_8246_out0;
assign v_RM_11368_out0 = v_S_8928_out0;
assign v_RM_11832_out0 = v_S_9392_out0;
assign v_G1_7783_out0 = ((v_RD_5928_out0 && !v_RM_11368_out0) || (!v_RD_5928_out0) && v_RM_11368_out0);
assign v_G1_8247_out0 = ((v_RD_6392_out0 && !v_RM_11832_out0) || (!v_RD_6392_out0) && v_RM_11832_out0);
assign v_G2_12319_out0 = v_RD_5928_out0 && v_RM_11368_out0;
assign v_G2_12783_out0 = v_RD_6392_out0 && v_RM_11832_out0;
assign v_CARRY_4928_out0 = v_G2_12319_out0;
assign v_CARRY_5392_out0 = v_G2_12783_out0;
assign v_S_8929_out0 = v_G1_7783_out0;
assign v_S_9393_out0 = v_G1_8247_out0;
assign v_S_1250_out0 = v_S_8929_out0;
assign v_S_1474_out0 = v_S_9393_out0;
assign v_G1_4026_out0 = v_CARRY_4928_out0 || v_CARRY_4927_out0;
assign v_G1_4250_out0 = v_CARRY_5392_out0 || v_CARRY_5391_out0;
assign v_COUT_718_out0 = v_G1_4026_out0;
assign v_COUT_942_out0 = v_G1_4250_out0;
assign v__10653_out0 = { v__4551_out0,v_S_1250_out0 };
assign v__10668_out0 = { v__4566_out0,v_S_1474_out0 };
assign v__10948_out0 = { v__10653_out0,v_COUT_718_out0 };
assign v__10963_out0 = { v__10668_out0,v_COUT_942_out0 };
assign v_COUT_10918_out0 = v__10948_out0;
assign v_COUT_10933_out0 = v__10963_out0;
assign v_CIN_2359_out0 = v_COUT_10918_out0;
assign v_CIN_2374_out0 = v_COUT_10933_out0;
assign v__472_out0 = v_CIN_2359_out0[8:8];
assign v__487_out0 = v_CIN_2374_out0[8:8];
assign v__1777_out0 = v_CIN_2359_out0[6:6];
assign v__1792_out0 = v_CIN_2374_out0[6:6];
assign v__2159_out0 = v_CIN_2359_out0[3:3];
assign v__2174_out0 = v_CIN_2374_out0[3:3];
assign v__2198_out0 = v_CIN_2359_out0[15:15];
assign v__2212_out0 = v_CIN_2374_out0[15:15];
assign v__2506_out0 = v_CIN_2359_out0[0:0];
assign v__2521_out0 = v_CIN_2374_out0[0:0];
assign v__3055_out0 = v_CIN_2359_out0[9:9];
assign v__3070_out0 = v_CIN_2374_out0[9:9];
assign v__3089_out0 = v_CIN_2359_out0[2:2];
assign v__3104_out0 = v_CIN_2374_out0[2:2];
assign v__3143_out0 = v_CIN_2359_out0[7:7];
assign v__3158_out0 = v_CIN_2374_out0[7:7];
assign v__3827_out0 = v_CIN_2359_out0[1:1];
assign v__3842_out0 = v_CIN_2374_out0[1:1];
assign v__3865_out0 = v_CIN_2359_out0[10:10];
assign v__3880_out0 = v_CIN_2374_out0[10:10];
assign v__6804_out0 = v_CIN_2359_out0[11:11];
assign v__6819_out0 = v_CIN_2374_out0[11:11];
assign v__7648_out0 = v_CIN_2359_out0[12:12];
assign v__7663_out0 = v_CIN_2374_out0[12:12];
assign v__8703_out0 = v_CIN_2359_out0[13:13];
assign v__8718_out0 = v_CIN_2374_out0[13:13];
assign v__8773_out0 = v_CIN_2359_out0[14:14];
assign v__8788_out0 = v_CIN_2374_out0[14:14];
assign v__10723_out0 = v_CIN_2359_out0[5:5];
assign v__10738_out0 = v_CIN_2374_out0[5:5];
assign v__13452_out0 = v_CIN_2359_out0[4:4];
assign v__13467_out0 = v_CIN_2374_out0[4:4];
assign v_RM_3414_out0 = v__7648_out0;
assign v_RM_3415_out0 = v__8773_out0;
assign v_RM_3417_out0 = v__10723_out0;
assign v_RM_3418_out0 = v__13452_out0;
assign v_RM_3419_out0 = v__8703_out0;
assign v_RM_3420_out0 = v__3055_out0;
assign v_RM_3421_out0 = v__3865_out0;
assign v_RM_3422_out0 = v__3827_out0;
assign v_RM_3423_out0 = v__2159_out0;
assign v_RM_3424_out0 = v__1777_out0;
assign v_RM_3425_out0 = v__3143_out0;
assign v_RM_3426_out0 = v__6804_out0;
assign v_RM_3427_out0 = v__472_out0;
assign v_RM_3428_out0 = v__3089_out0;
assign v_RM_3638_out0 = v__7663_out0;
assign v_RM_3639_out0 = v__8788_out0;
assign v_RM_3641_out0 = v__10738_out0;
assign v_RM_3642_out0 = v__13467_out0;
assign v_RM_3643_out0 = v__8718_out0;
assign v_RM_3644_out0 = v__3070_out0;
assign v_RM_3645_out0 = v__3880_out0;
assign v_RM_3646_out0 = v__3842_out0;
assign v_RM_3647_out0 = v__2174_out0;
assign v_RM_3648_out0 = v__1792_out0;
assign v_RM_3649_out0 = v__3158_out0;
assign v_RM_3650_out0 = v__6819_out0;
assign v_RM_3651_out0 = v__487_out0;
assign v_RM_3652_out0 = v__3104_out0;
assign v_CIN_9869_out0 = v__2198_out0;
assign v_CIN_10093_out0 = v__2212_out0;
assign v_RM_11437_out0 = v__2506_out0;
assign v_RM_11901_out0 = v__2521_out0;
assign v_RD_5990_out0 = v_CIN_9869_out0;
assign v_RD_6454_out0 = v_CIN_10093_out0;
assign v_G1_7852_out0 = ((v_RD_5997_out0 && !v_RM_11437_out0) || (!v_RD_5997_out0) && v_RM_11437_out0);
assign v_G1_8316_out0 = ((v_RD_6461_out0 && !v_RM_11901_out0) || (!v_RD_6461_out0) && v_RM_11901_out0);
assign v_RM_11425_out0 = v_RM_3414_out0;
assign v_RM_11427_out0 = v_RM_3415_out0;
assign v_RM_11431_out0 = v_RM_3417_out0;
assign v_RM_11433_out0 = v_RM_3418_out0;
assign v_RM_11435_out0 = v_RM_3419_out0;
assign v_RM_11438_out0 = v_RM_3420_out0;
assign v_RM_11440_out0 = v_RM_3421_out0;
assign v_RM_11442_out0 = v_RM_3422_out0;
assign v_RM_11444_out0 = v_RM_3423_out0;
assign v_RM_11446_out0 = v_RM_3424_out0;
assign v_RM_11448_out0 = v_RM_3425_out0;
assign v_RM_11450_out0 = v_RM_3426_out0;
assign v_RM_11452_out0 = v_RM_3427_out0;
assign v_RM_11454_out0 = v_RM_3428_out0;
assign v_RM_11889_out0 = v_RM_3638_out0;
assign v_RM_11891_out0 = v_RM_3639_out0;
assign v_RM_11895_out0 = v_RM_3641_out0;
assign v_RM_11897_out0 = v_RM_3642_out0;
assign v_RM_11899_out0 = v_RM_3643_out0;
assign v_RM_11902_out0 = v_RM_3644_out0;
assign v_RM_11904_out0 = v_RM_3645_out0;
assign v_RM_11906_out0 = v_RM_3646_out0;
assign v_RM_11908_out0 = v_RM_3647_out0;
assign v_RM_11910_out0 = v_RM_3648_out0;
assign v_RM_11912_out0 = v_RM_3649_out0;
assign v_RM_11914_out0 = v_RM_3650_out0;
assign v_RM_11916_out0 = v_RM_3651_out0;
assign v_RM_11918_out0 = v_RM_3652_out0;
assign v_G2_12388_out0 = v_RD_5997_out0 && v_RM_11437_out0;
assign v_G2_12852_out0 = v_RD_6461_out0 && v_RM_11901_out0;
assign v_CARRY_4997_out0 = v_G2_12388_out0;
assign v_CARRY_5461_out0 = v_G2_12852_out0;
assign v_G1_7840_out0 = ((v_RD_5985_out0 && !v_RM_11425_out0) || (!v_RD_5985_out0) && v_RM_11425_out0);
assign v_G1_7842_out0 = ((v_RD_5987_out0 && !v_RM_11427_out0) || (!v_RD_5987_out0) && v_RM_11427_out0);
assign v_G1_7846_out0 = ((v_RD_5991_out0 && !v_RM_11431_out0) || (!v_RD_5991_out0) && v_RM_11431_out0);
assign v_G1_7848_out0 = ((v_RD_5993_out0 && !v_RM_11433_out0) || (!v_RD_5993_out0) && v_RM_11433_out0);
assign v_G1_7850_out0 = ((v_RD_5995_out0 && !v_RM_11435_out0) || (!v_RD_5995_out0) && v_RM_11435_out0);
assign v_G1_7853_out0 = ((v_RD_5998_out0 && !v_RM_11438_out0) || (!v_RD_5998_out0) && v_RM_11438_out0);
assign v_G1_7855_out0 = ((v_RD_6000_out0 && !v_RM_11440_out0) || (!v_RD_6000_out0) && v_RM_11440_out0);
assign v_G1_7857_out0 = ((v_RD_6002_out0 && !v_RM_11442_out0) || (!v_RD_6002_out0) && v_RM_11442_out0);
assign v_G1_7859_out0 = ((v_RD_6004_out0 && !v_RM_11444_out0) || (!v_RD_6004_out0) && v_RM_11444_out0);
assign v_G1_7861_out0 = ((v_RD_6006_out0 && !v_RM_11446_out0) || (!v_RD_6006_out0) && v_RM_11446_out0);
assign v_G1_7863_out0 = ((v_RD_6008_out0 && !v_RM_11448_out0) || (!v_RD_6008_out0) && v_RM_11448_out0);
assign v_G1_7865_out0 = ((v_RD_6010_out0 && !v_RM_11450_out0) || (!v_RD_6010_out0) && v_RM_11450_out0);
assign v_G1_7867_out0 = ((v_RD_6012_out0 && !v_RM_11452_out0) || (!v_RD_6012_out0) && v_RM_11452_out0);
assign v_G1_7869_out0 = ((v_RD_6014_out0 && !v_RM_11454_out0) || (!v_RD_6014_out0) && v_RM_11454_out0);
assign v_G1_8304_out0 = ((v_RD_6449_out0 && !v_RM_11889_out0) || (!v_RD_6449_out0) && v_RM_11889_out0);
assign v_G1_8306_out0 = ((v_RD_6451_out0 && !v_RM_11891_out0) || (!v_RD_6451_out0) && v_RM_11891_out0);
assign v_G1_8310_out0 = ((v_RD_6455_out0 && !v_RM_11895_out0) || (!v_RD_6455_out0) && v_RM_11895_out0);
assign v_G1_8312_out0 = ((v_RD_6457_out0 && !v_RM_11897_out0) || (!v_RD_6457_out0) && v_RM_11897_out0);
assign v_G1_8314_out0 = ((v_RD_6459_out0 && !v_RM_11899_out0) || (!v_RD_6459_out0) && v_RM_11899_out0);
assign v_G1_8317_out0 = ((v_RD_6462_out0 && !v_RM_11902_out0) || (!v_RD_6462_out0) && v_RM_11902_out0);
assign v_G1_8319_out0 = ((v_RD_6464_out0 && !v_RM_11904_out0) || (!v_RD_6464_out0) && v_RM_11904_out0);
assign v_G1_8321_out0 = ((v_RD_6466_out0 && !v_RM_11906_out0) || (!v_RD_6466_out0) && v_RM_11906_out0);
assign v_G1_8323_out0 = ((v_RD_6468_out0 && !v_RM_11908_out0) || (!v_RD_6468_out0) && v_RM_11908_out0);
assign v_G1_8325_out0 = ((v_RD_6470_out0 && !v_RM_11910_out0) || (!v_RD_6470_out0) && v_RM_11910_out0);
assign v_G1_8327_out0 = ((v_RD_6472_out0 && !v_RM_11912_out0) || (!v_RD_6472_out0) && v_RM_11912_out0);
assign v_G1_8329_out0 = ((v_RD_6474_out0 && !v_RM_11914_out0) || (!v_RD_6474_out0) && v_RM_11914_out0);
assign v_G1_8331_out0 = ((v_RD_6476_out0 && !v_RM_11916_out0) || (!v_RD_6476_out0) && v_RM_11916_out0);
assign v_G1_8333_out0 = ((v_RD_6478_out0 && !v_RM_11918_out0) || (!v_RD_6478_out0) && v_RM_11918_out0);
assign v_S_8998_out0 = v_G1_7852_out0;
assign v_S_9462_out0 = v_G1_8316_out0;
assign v_G2_12376_out0 = v_RD_5985_out0 && v_RM_11425_out0;
assign v_G2_12378_out0 = v_RD_5987_out0 && v_RM_11427_out0;
assign v_G2_12382_out0 = v_RD_5991_out0 && v_RM_11431_out0;
assign v_G2_12384_out0 = v_RD_5993_out0 && v_RM_11433_out0;
assign v_G2_12386_out0 = v_RD_5995_out0 && v_RM_11435_out0;
assign v_G2_12389_out0 = v_RD_5998_out0 && v_RM_11438_out0;
assign v_G2_12391_out0 = v_RD_6000_out0 && v_RM_11440_out0;
assign v_G2_12393_out0 = v_RD_6002_out0 && v_RM_11442_out0;
assign v_G2_12395_out0 = v_RD_6004_out0 && v_RM_11444_out0;
assign v_G2_12397_out0 = v_RD_6006_out0 && v_RM_11446_out0;
assign v_G2_12399_out0 = v_RD_6008_out0 && v_RM_11448_out0;
assign v_G2_12401_out0 = v_RD_6010_out0 && v_RM_11450_out0;
assign v_G2_12403_out0 = v_RD_6012_out0 && v_RM_11452_out0;
assign v_G2_12405_out0 = v_RD_6014_out0 && v_RM_11454_out0;
assign v_G2_12840_out0 = v_RD_6449_out0 && v_RM_11889_out0;
assign v_G2_12842_out0 = v_RD_6451_out0 && v_RM_11891_out0;
assign v_G2_12846_out0 = v_RD_6455_out0 && v_RM_11895_out0;
assign v_G2_12848_out0 = v_RD_6457_out0 && v_RM_11897_out0;
assign v_G2_12850_out0 = v_RD_6459_out0 && v_RM_11899_out0;
assign v_G2_12853_out0 = v_RD_6462_out0 && v_RM_11902_out0;
assign v_G2_12855_out0 = v_RD_6464_out0 && v_RM_11904_out0;
assign v_G2_12857_out0 = v_RD_6466_out0 && v_RM_11906_out0;
assign v_G2_12859_out0 = v_RD_6468_out0 && v_RM_11908_out0;
assign v_G2_12861_out0 = v_RD_6470_out0 && v_RM_11910_out0;
assign v_G2_12863_out0 = v_RD_6472_out0 && v_RM_11912_out0;
assign v_G2_12865_out0 = v_RD_6474_out0 && v_RM_11914_out0;
assign v_G2_12867_out0 = v_RD_6476_out0 && v_RM_11916_out0;
assign v_G2_12869_out0 = v_RD_6478_out0 && v_RM_11918_out0;
assign v_S_4669_out0 = v_S_8998_out0;
assign v_S_4684_out0 = v_S_9462_out0;
assign v_CARRY_4985_out0 = v_G2_12376_out0;
assign v_CARRY_4987_out0 = v_G2_12378_out0;
assign v_CARRY_4991_out0 = v_G2_12382_out0;
assign v_CARRY_4993_out0 = v_G2_12384_out0;
assign v_CARRY_4995_out0 = v_G2_12386_out0;
assign v_CARRY_4998_out0 = v_G2_12389_out0;
assign v_CARRY_5000_out0 = v_G2_12391_out0;
assign v_CARRY_5002_out0 = v_G2_12393_out0;
assign v_CARRY_5004_out0 = v_G2_12395_out0;
assign v_CARRY_5006_out0 = v_G2_12397_out0;
assign v_CARRY_5008_out0 = v_G2_12399_out0;
assign v_CARRY_5010_out0 = v_G2_12401_out0;
assign v_CARRY_5012_out0 = v_G2_12403_out0;
assign v_CARRY_5014_out0 = v_G2_12405_out0;
assign v_CARRY_5449_out0 = v_G2_12840_out0;
assign v_CARRY_5451_out0 = v_G2_12842_out0;
assign v_CARRY_5455_out0 = v_G2_12846_out0;
assign v_CARRY_5457_out0 = v_G2_12848_out0;
assign v_CARRY_5459_out0 = v_G2_12850_out0;
assign v_CARRY_5462_out0 = v_G2_12853_out0;
assign v_CARRY_5464_out0 = v_G2_12855_out0;
assign v_CARRY_5466_out0 = v_G2_12857_out0;
assign v_CARRY_5468_out0 = v_G2_12859_out0;
assign v_CARRY_5470_out0 = v_G2_12861_out0;
assign v_CARRY_5472_out0 = v_G2_12863_out0;
assign v_CARRY_5474_out0 = v_G2_12865_out0;
assign v_CARRY_5476_out0 = v_G2_12867_out0;
assign v_CARRY_5478_out0 = v_G2_12869_out0;
assign v_S_8986_out0 = v_G1_7840_out0;
assign v_S_8988_out0 = v_G1_7842_out0;
assign v_S_8992_out0 = v_G1_7846_out0;
assign v_S_8994_out0 = v_G1_7848_out0;
assign v_S_8996_out0 = v_G1_7850_out0;
assign v_S_8999_out0 = v_G1_7853_out0;
assign v_S_9001_out0 = v_G1_7855_out0;
assign v_S_9003_out0 = v_G1_7857_out0;
assign v_S_9005_out0 = v_G1_7859_out0;
assign v_S_9007_out0 = v_G1_7861_out0;
assign v_S_9009_out0 = v_G1_7863_out0;
assign v_S_9011_out0 = v_G1_7865_out0;
assign v_S_9013_out0 = v_G1_7867_out0;
assign v_S_9015_out0 = v_G1_7869_out0;
assign v_S_9450_out0 = v_G1_8304_out0;
assign v_S_9452_out0 = v_G1_8306_out0;
assign v_S_9456_out0 = v_G1_8310_out0;
assign v_S_9458_out0 = v_G1_8312_out0;
assign v_S_9460_out0 = v_G1_8314_out0;
assign v_S_9463_out0 = v_G1_8317_out0;
assign v_S_9465_out0 = v_G1_8319_out0;
assign v_S_9467_out0 = v_G1_8321_out0;
assign v_S_9469_out0 = v_G1_8323_out0;
assign v_S_9471_out0 = v_G1_8325_out0;
assign v_S_9473_out0 = v_G1_8327_out0;
assign v_S_9475_out0 = v_G1_8329_out0;
assign v_S_9477_out0 = v_G1_8331_out0;
assign v_S_9479_out0 = v_G1_8333_out0;
assign v_CIN_9875_out0 = v_CARRY_4997_out0;
assign v_CIN_10099_out0 = v_CARRY_5461_out0;
assign v__4529_out0 = { v__1716_out0,v_S_4669_out0 };
assign v__4530_out0 = { v__1717_out0,v_S_4684_out0 };
assign v_RD_6003_out0 = v_CIN_9875_out0;
assign v_RD_6467_out0 = v_CIN_10099_out0;
assign v_RM_11426_out0 = v_S_8986_out0;
assign v_RM_11428_out0 = v_S_8988_out0;
assign v_RM_11432_out0 = v_S_8992_out0;
assign v_RM_11434_out0 = v_S_8994_out0;
assign v_RM_11436_out0 = v_S_8996_out0;
assign v_RM_11439_out0 = v_S_8999_out0;
assign v_RM_11441_out0 = v_S_9001_out0;
assign v_RM_11443_out0 = v_S_9003_out0;
assign v_RM_11445_out0 = v_S_9005_out0;
assign v_RM_11447_out0 = v_S_9007_out0;
assign v_RM_11449_out0 = v_S_9009_out0;
assign v_RM_11451_out0 = v_S_9011_out0;
assign v_RM_11453_out0 = v_S_9013_out0;
assign v_RM_11455_out0 = v_S_9015_out0;
assign v_RM_11890_out0 = v_S_9450_out0;
assign v_RM_11892_out0 = v_S_9452_out0;
assign v_RM_11896_out0 = v_S_9456_out0;
assign v_RM_11898_out0 = v_S_9458_out0;
assign v_RM_11900_out0 = v_S_9460_out0;
assign v_RM_11903_out0 = v_S_9463_out0;
assign v_RM_11905_out0 = v_S_9465_out0;
assign v_RM_11907_out0 = v_S_9467_out0;
assign v_RM_11909_out0 = v_S_9469_out0;
assign v_RM_11911_out0 = v_S_9471_out0;
assign v_RM_11913_out0 = v_S_9473_out0;
assign v_RM_11915_out0 = v_S_9475_out0;
assign v_RM_11917_out0 = v_S_9477_out0;
assign v_RM_11919_out0 = v_S_9479_out0;
assign v_G1_7858_out0 = ((v_RD_6003_out0 && !v_RM_11443_out0) || (!v_RD_6003_out0) && v_RM_11443_out0);
assign v_G1_8322_out0 = ((v_RD_6467_out0 && !v_RM_11907_out0) || (!v_RD_6467_out0) && v_RM_11907_out0);
assign v_G2_12394_out0 = v_RD_6003_out0 && v_RM_11443_out0;
assign v_G2_12858_out0 = v_RD_6467_out0 && v_RM_11907_out0;
assign v_CARRY_5003_out0 = v_G2_12394_out0;
assign v_CARRY_5467_out0 = v_G2_12858_out0;
assign v_S_9004_out0 = v_G1_7858_out0;
assign v_S_9468_out0 = v_G1_8322_out0;
assign v_S_1286_out0 = v_S_9004_out0;
assign v_S_1510_out0 = v_S_9468_out0;
assign v_G1_4062_out0 = v_CARRY_5003_out0 || v_CARRY_5002_out0;
assign v_G1_4286_out0 = v_CARRY_5467_out0 || v_CARRY_5466_out0;
assign v_COUT_754_out0 = v_G1_4062_out0;
assign v_COUT_978_out0 = v_G1_4286_out0;
assign v_CIN_9881_out0 = v_COUT_754_out0;
assign v_CIN_10105_out0 = v_COUT_978_out0;
assign v_RD_6015_out0 = v_CIN_9881_out0;
assign v_RD_6479_out0 = v_CIN_10105_out0;
assign v_G1_7870_out0 = ((v_RD_6015_out0 && !v_RM_11455_out0) || (!v_RD_6015_out0) && v_RM_11455_out0);
assign v_G1_8334_out0 = ((v_RD_6479_out0 && !v_RM_11919_out0) || (!v_RD_6479_out0) && v_RM_11919_out0);
assign v_G2_12406_out0 = v_RD_6015_out0 && v_RM_11455_out0;
assign v_G2_12870_out0 = v_RD_6479_out0 && v_RM_11919_out0;
assign v_CARRY_5015_out0 = v_G2_12406_out0;
assign v_CARRY_5479_out0 = v_G2_12870_out0;
assign v_S_9016_out0 = v_G1_7870_out0;
assign v_S_9480_out0 = v_G1_8334_out0;
assign v_S_1292_out0 = v_S_9016_out0;
assign v_S_1516_out0 = v_S_9480_out0;
assign v_G1_4068_out0 = v_CARRY_5015_out0 || v_CARRY_5014_out0;
assign v_G1_4292_out0 = v_CARRY_5479_out0 || v_CARRY_5478_out0;
assign v_COUT_760_out0 = v_G1_4068_out0;
assign v_COUT_984_out0 = v_G1_4292_out0;
assign v__4786_out0 = { v_S_1286_out0,v_S_1292_out0 };
assign v__4801_out0 = { v_S_1510_out0,v_S_1516_out0 };
assign v_CIN_9876_out0 = v_COUT_760_out0;
assign v_CIN_10100_out0 = v_COUT_984_out0;
assign v_RD_6005_out0 = v_CIN_9876_out0;
assign v_RD_6469_out0 = v_CIN_10100_out0;
assign v_G1_7860_out0 = ((v_RD_6005_out0 && !v_RM_11445_out0) || (!v_RD_6005_out0) && v_RM_11445_out0);
assign v_G1_8324_out0 = ((v_RD_6469_out0 && !v_RM_11909_out0) || (!v_RD_6469_out0) && v_RM_11909_out0);
assign v_G2_12396_out0 = v_RD_6005_out0 && v_RM_11445_out0;
assign v_G2_12860_out0 = v_RD_6469_out0 && v_RM_11909_out0;
assign v_CARRY_5005_out0 = v_G2_12396_out0;
assign v_CARRY_5469_out0 = v_G2_12860_out0;
assign v_S_9006_out0 = v_G1_7860_out0;
assign v_S_9470_out0 = v_G1_8324_out0;
assign v_S_1287_out0 = v_S_9006_out0;
assign v_S_1511_out0 = v_S_9470_out0;
assign v_G1_4063_out0 = v_CARRY_5005_out0 || v_CARRY_5004_out0;
assign v_G1_4287_out0 = v_CARRY_5469_out0 || v_CARRY_5468_out0;
assign v_COUT_755_out0 = v_G1_4063_out0;
assign v_COUT_979_out0 = v_G1_4287_out0;
assign v__2556_out0 = { v__4786_out0,v_S_1287_out0 };
assign v__2571_out0 = { v__4801_out0,v_S_1511_out0 };
assign v_CIN_9871_out0 = v_COUT_755_out0;
assign v_CIN_10095_out0 = v_COUT_979_out0;
assign v_RD_5994_out0 = v_CIN_9871_out0;
assign v_RD_6458_out0 = v_CIN_10095_out0;
assign v_G1_7849_out0 = ((v_RD_5994_out0 && !v_RM_11434_out0) || (!v_RD_5994_out0) && v_RM_11434_out0);
assign v_G1_8313_out0 = ((v_RD_6458_out0 && !v_RM_11898_out0) || (!v_RD_6458_out0) && v_RM_11898_out0);
assign v_G2_12385_out0 = v_RD_5994_out0 && v_RM_11434_out0;
assign v_G2_12849_out0 = v_RD_6458_out0 && v_RM_11898_out0;
assign v_CARRY_4994_out0 = v_G2_12385_out0;
assign v_CARRY_5458_out0 = v_G2_12849_out0;
assign v_S_8995_out0 = v_G1_7849_out0;
assign v_S_9459_out0 = v_G1_8313_out0;
assign v_S_1282_out0 = v_S_8995_out0;
assign v_S_1506_out0 = v_S_9459_out0;
assign v_G1_4058_out0 = v_CARRY_4994_out0 || v_CARRY_4993_out0;
assign v_G1_4282_out0 = v_CARRY_5458_out0 || v_CARRY_5457_out0;
assign v_COUT_750_out0 = v_G1_4058_out0;
assign v_COUT_974_out0 = v_G1_4282_out0;
assign v__7036_out0 = { v__2556_out0,v_S_1282_out0 };
assign v__7051_out0 = { v__2571_out0,v_S_1506_out0 };
assign v_CIN_9870_out0 = v_COUT_750_out0;
assign v_CIN_10094_out0 = v_COUT_974_out0;
assign v_RD_5992_out0 = v_CIN_9870_out0;
assign v_RD_6456_out0 = v_CIN_10094_out0;
assign v_G1_7847_out0 = ((v_RD_5992_out0 && !v_RM_11432_out0) || (!v_RD_5992_out0) && v_RM_11432_out0);
assign v_G1_8311_out0 = ((v_RD_6456_out0 && !v_RM_11896_out0) || (!v_RD_6456_out0) && v_RM_11896_out0);
assign v_G2_12383_out0 = v_RD_5992_out0 && v_RM_11432_out0;
assign v_G2_12847_out0 = v_RD_6456_out0 && v_RM_11896_out0;
assign v_CARRY_4992_out0 = v_G2_12383_out0;
assign v_CARRY_5456_out0 = v_G2_12847_out0;
assign v_S_8993_out0 = v_G1_7847_out0;
assign v_S_9457_out0 = v_G1_8311_out0;
assign v_S_1281_out0 = v_S_8993_out0;
assign v_S_1505_out0 = v_S_9457_out0;
assign v_G1_4057_out0 = v_CARRY_4992_out0 || v_CARRY_4991_out0;
assign v_G1_4281_out0 = v_CARRY_5456_out0 || v_CARRY_5455_out0;
assign v_COUT_749_out0 = v_G1_4057_out0;
assign v_COUT_973_out0 = v_G1_4281_out0;
assign v__13522_out0 = { v__7036_out0,v_S_1281_out0 };
assign v__13537_out0 = { v__7051_out0,v_S_1505_out0 };
assign v_CIN_9877_out0 = v_COUT_749_out0;
assign v_CIN_10101_out0 = v_COUT_973_out0;
assign v_RD_6007_out0 = v_CIN_9877_out0;
assign v_RD_6471_out0 = v_CIN_10101_out0;
assign v_G1_7862_out0 = ((v_RD_6007_out0 && !v_RM_11447_out0) || (!v_RD_6007_out0) && v_RM_11447_out0);
assign v_G1_8326_out0 = ((v_RD_6471_out0 && !v_RM_11911_out0) || (!v_RD_6471_out0) && v_RM_11911_out0);
assign v_G2_12398_out0 = v_RD_6007_out0 && v_RM_11447_out0;
assign v_G2_12862_out0 = v_RD_6471_out0 && v_RM_11911_out0;
assign v_CARRY_5007_out0 = v_G2_12398_out0;
assign v_CARRY_5471_out0 = v_G2_12862_out0;
assign v_S_9008_out0 = v_G1_7862_out0;
assign v_S_9472_out0 = v_G1_8326_out0;
assign v_S_1288_out0 = v_S_9008_out0;
assign v_S_1512_out0 = v_S_9472_out0;
assign v_G1_4064_out0 = v_CARRY_5007_out0 || v_CARRY_5006_out0;
assign v_G1_4288_out0 = v_CARRY_5471_out0 || v_CARRY_5470_out0;
assign v_COUT_756_out0 = v_G1_4064_out0;
assign v_COUT_980_out0 = v_G1_4288_out0;
assign v__3315_out0 = { v__13522_out0,v_S_1288_out0 };
assign v__3330_out0 = { v__13537_out0,v_S_1512_out0 };
assign v_CIN_9878_out0 = v_COUT_756_out0;
assign v_CIN_10102_out0 = v_COUT_980_out0;
assign v_RD_6009_out0 = v_CIN_9878_out0;
assign v_RD_6473_out0 = v_CIN_10102_out0;
assign v_G1_7864_out0 = ((v_RD_6009_out0 && !v_RM_11449_out0) || (!v_RD_6009_out0) && v_RM_11449_out0);
assign v_G1_8328_out0 = ((v_RD_6473_out0 && !v_RM_11913_out0) || (!v_RD_6473_out0) && v_RM_11913_out0);
assign v_G2_12400_out0 = v_RD_6009_out0 && v_RM_11449_out0;
assign v_G2_12864_out0 = v_RD_6473_out0 && v_RM_11913_out0;
assign v_CARRY_5009_out0 = v_G2_12400_out0;
assign v_CARRY_5473_out0 = v_G2_12864_out0;
assign v_S_9010_out0 = v_G1_7864_out0;
assign v_S_9474_out0 = v_G1_8328_out0;
assign v_S_1289_out0 = v_S_9010_out0;
assign v_S_1513_out0 = v_S_9474_out0;
assign v_G1_4065_out0 = v_CARRY_5009_out0 || v_CARRY_5008_out0;
assign v_G1_4289_out0 = v_CARRY_5473_out0 || v_CARRY_5472_out0;
assign v_COUT_757_out0 = v_G1_4065_out0;
assign v_COUT_981_out0 = v_G1_4289_out0;
assign v__7151_out0 = { v__3315_out0,v_S_1289_out0 };
assign v__7166_out0 = { v__3330_out0,v_S_1513_out0 };
assign v_CIN_9880_out0 = v_COUT_757_out0;
assign v_CIN_10104_out0 = v_COUT_981_out0;
assign v_RD_6013_out0 = v_CIN_9880_out0;
assign v_RD_6477_out0 = v_CIN_10104_out0;
assign v_G1_7868_out0 = ((v_RD_6013_out0 && !v_RM_11453_out0) || (!v_RD_6013_out0) && v_RM_11453_out0);
assign v_G1_8332_out0 = ((v_RD_6477_out0 && !v_RM_11917_out0) || (!v_RD_6477_out0) && v_RM_11917_out0);
assign v_G2_12404_out0 = v_RD_6013_out0 && v_RM_11453_out0;
assign v_G2_12868_out0 = v_RD_6477_out0 && v_RM_11917_out0;
assign v_CARRY_5013_out0 = v_G2_12404_out0;
assign v_CARRY_5477_out0 = v_G2_12868_out0;
assign v_S_9014_out0 = v_G1_7868_out0;
assign v_S_9478_out0 = v_G1_8332_out0;
assign v_S_1291_out0 = v_S_9014_out0;
assign v_S_1515_out0 = v_S_9478_out0;
assign v_G1_4067_out0 = v_CARRY_5013_out0 || v_CARRY_5012_out0;
assign v_G1_4291_out0 = v_CARRY_5477_out0 || v_CARRY_5476_out0;
assign v_COUT_759_out0 = v_G1_4067_out0;
assign v_COUT_983_out0 = v_G1_4291_out0;
assign v__4753_out0 = { v__7151_out0,v_S_1291_out0 };
assign v__4768_out0 = { v__7166_out0,v_S_1515_out0 };
assign v_CIN_9873_out0 = v_COUT_759_out0;
assign v_CIN_10097_out0 = v_COUT_983_out0;
assign v_RD_5999_out0 = v_CIN_9873_out0;
assign v_RD_6463_out0 = v_CIN_10097_out0;
assign v_G1_7854_out0 = ((v_RD_5999_out0 && !v_RM_11439_out0) || (!v_RD_5999_out0) && v_RM_11439_out0);
assign v_G1_8318_out0 = ((v_RD_6463_out0 && !v_RM_11903_out0) || (!v_RD_6463_out0) && v_RM_11903_out0);
assign v_G2_12390_out0 = v_RD_5999_out0 && v_RM_11439_out0;
assign v_G2_12854_out0 = v_RD_6463_out0 && v_RM_11903_out0;
assign v_CARRY_4999_out0 = v_G2_12390_out0;
assign v_CARRY_5463_out0 = v_G2_12854_out0;
assign v_S_9000_out0 = v_G1_7854_out0;
assign v_S_9464_out0 = v_G1_8318_out0;
assign v_S_1284_out0 = v_S_9000_out0;
assign v_S_1508_out0 = v_S_9464_out0;
assign v_G1_4060_out0 = v_CARRY_4999_out0 || v_CARRY_4998_out0;
assign v_G1_4284_out0 = v_CARRY_5463_out0 || v_CARRY_5462_out0;
assign v_COUT_752_out0 = v_G1_4060_out0;
assign v_COUT_976_out0 = v_G1_4284_out0;
assign v__6930_out0 = { v__4753_out0,v_S_1284_out0 };
assign v__6945_out0 = { v__4768_out0,v_S_1508_out0 };
assign v_CIN_9874_out0 = v_COUT_752_out0;
assign v_CIN_10098_out0 = v_COUT_976_out0;
assign v_RD_6001_out0 = v_CIN_9874_out0;
assign v_RD_6465_out0 = v_CIN_10098_out0;
assign v_G1_7856_out0 = ((v_RD_6001_out0 && !v_RM_11441_out0) || (!v_RD_6001_out0) && v_RM_11441_out0);
assign v_G1_8320_out0 = ((v_RD_6465_out0 && !v_RM_11905_out0) || (!v_RD_6465_out0) && v_RM_11905_out0);
assign v_G2_12392_out0 = v_RD_6001_out0 && v_RM_11441_out0;
assign v_G2_12856_out0 = v_RD_6465_out0 && v_RM_11905_out0;
assign v_CARRY_5001_out0 = v_G2_12392_out0;
assign v_CARRY_5465_out0 = v_G2_12856_out0;
assign v_S_9002_out0 = v_G1_7856_out0;
assign v_S_9466_out0 = v_G1_8320_out0;
assign v_S_1285_out0 = v_S_9002_out0;
assign v_S_1509_out0 = v_S_9466_out0;
assign v_G1_4061_out0 = v_CARRY_5001_out0 || v_CARRY_5000_out0;
assign v_G1_4285_out0 = v_CARRY_5465_out0 || v_CARRY_5464_out0;
assign v_COUT_753_out0 = v_G1_4061_out0;
assign v_COUT_977_out0 = v_G1_4285_out0;
assign v__5806_out0 = { v__6930_out0,v_S_1285_out0 };
assign v__5821_out0 = { v__6945_out0,v_S_1509_out0 };
assign v_CIN_9879_out0 = v_COUT_753_out0;
assign v_CIN_10103_out0 = v_COUT_977_out0;
assign v_RD_6011_out0 = v_CIN_9879_out0;
assign v_RD_6475_out0 = v_CIN_10103_out0;
assign v_G1_7866_out0 = ((v_RD_6011_out0 && !v_RM_11451_out0) || (!v_RD_6011_out0) && v_RM_11451_out0);
assign v_G1_8330_out0 = ((v_RD_6475_out0 && !v_RM_11915_out0) || (!v_RD_6475_out0) && v_RM_11915_out0);
assign v_G2_12402_out0 = v_RD_6011_out0 && v_RM_11451_out0;
assign v_G2_12866_out0 = v_RD_6475_out0 && v_RM_11915_out0;
assign v_CARRY_5011_out0 = v_G2_12402_out0;
assign v_CARRY_5475_out0 = v_G2_12866_out0;
assign v_S_9012_out0 = v_G1_7866_out0;
assign v_S_9476_out0 = v_G1_8330_out0;
assign v_S_1290_out0 = v_S_9012_out0;
assign v_S_1514_out0 = v_S_9476_out0;
assign v_G1_4066_out0 = v_CARRY_5011_out0 || v_CARRY_5010_out0;
assign v_G1_4290_out0 = v_CARRY_5475_out0 || v_CARRY_5474_out0;
assign v_COUT_758_out0 = v_G1_4066_out0;
assign v_COUT_982_out0 = v_G1_4290_out0;
assign v__2030_out0 = { v__5806_out0,v_S_1290_out0 };
assign v__2045_out0 = { v__5821_out0,v_S_1514_out0 };
assign v_CIN_9867_out0 = v_COUT_758_out0;
assign v_CIN_10091_out0 = v_COUT_982_out0;
assign v_RD_5986_out0 = v_CIN_9867_out0;
assign v_RD_6450_out0 = v_CIN_10091_out0;
assign v_G1_7841_out0 = ((v_RD_5986_out0 && !v_RM_11426_out0) || (!v_RD_5986_out0) && v_RM_11426_out0);
assign v_G1_8305_out0 = ((v_RD_6450_out0 && !v_RM_11890_out0) || (!v_RD_6450_out0) && v_RM_11890_out0);
assign v_G2_12377_out0 = v_RD_5986_out0 && v_RM_11426_out0;
assign v_G2_12841_out0 = v_RD_6450_out0 && v_RM_11890_out0;
assign v_CARRY_4986_out0 = v_G2_12377_out0;
assign v_CARRY_5450_out0 = v_G2_12841_out0;
assign v_S_8987_out0 = v_G1_7841_out0;
assign v_S_9451_out0 = v_G1_8305_out0;
assign v_S_1278_out0 = v_S_8987_out0;
assign v_S_1502_out0 = v_S_9451_out0;
assign v_G1_4054_out0 = v_CARRY_4986_out0 || v_CARRY_4985_out0;
assign v_G1_4278_out0 = v_CARRY_5450_out0 || v_CARRY_5449_out0;
assign v_COUT_746_out0 = v_G1_4054_out0;
assign v_COUT_970_out0 = v_G1_4278_out0;
assign v__2797_out0 = { v__2030_out0,v_S_1278_out0 };
assign v__2812_out0 = { v__2045_out0,v_S_1502_out0 };
assign v_CIN_9872_out0 = v_COUT_746_out0;
assign v_CIN_10096_out0 = v_COUT_970_out0;
assign v_RD_5996_out0 = v_CIN_9872_out0;
assign v_RD_6460_out0 = v_CIN_10096_out0;
assign v_G1_7851_out0 = ((v_RD_5996_out0 && !v_RM_11436_out0) || (!v_RD_5996_out0) && v_RM_11436_out0);
assign v_G1_8315_out0 = ((v_RD_6460_out0 && !v_RM_11900_out0) || (!v_RD_6460_out0) && v_RM_11900_out0);
assign v_G2_12387_out0 = v_RD_5996_out0 && v_RM_11436_out0;
assign v_G2_12851_out0 = v_RD_6460_out0 && v_RM_11900_out0;
assign v_CARRY_4996_out0 = v_G2_12387_out0;
assign v_CARRY_5460_out0 = v_G2_12851_out0;
assign v_S_8997_out0 = v_G1_7851_out0;
assign v_S_9461_out0 = v_G1_8315_out0;
assign v_S_1283_out0 = v_S_8997_out0;
assign v_S_1507_out0 = v_S_9461_out0;
assign v_G1_4059_out0 = v_CARRY_4996_out0 || v_CARRY_4995_out0;
assign v_G1_4283_out0 = v_CARRY_5460_out0 || v_CARRY_5459_out0;
assign v_COUT_751_out0 = v_G1_4059_out0;
assign v_COUT_975_out0 = v_G1_4283_out0;
assign v__1829_out0 = { v__2797_out0,v_S_1283_out0 };
assign v__1844_out0 = { v__2812_out0,v_S_1507_out0 };
assign v_CIN_9868_out0 = v_COUT_751_out0;
assign v_CIN_10092_out0 = v_COUT_975_out0;
assign v_RD_5988_out0 = v_CIN_9868_out0;
assign v_RD_6452_out0 = v_CIN_10092_out0;
assign v_G1_7843_out0 = ((v_RD_5988_out0 && !v_RM_11428_out0) || (!v_RD_5988_out0) && v_RM_11428_out0);
assign v_G1_8307_out0 = ((v_RD_6452_out0 && !v_RM_11892_out0) || (!v_RD_6452_out0) && v_RM_11892_out0);
assign v_G2_12379_out0 = v_RD_5988_out0 && v_RM_11428_out0;
assign v_G2_12843_out0 = v_RD_6452_out0 && v_RM_11892_out0;
assign v_CARRY_4988_out0 = v_G2_12379_out0;
assign v_CARRY_5452_out0 = v_G2_12843_out0;
assign v_S_8989_out0 = v_G1_7843_out0;
assign v_S_9453_out0 = v_G1_8307_out0;
assign v_S_1279_out0 = v_S_8989_out0;
assign v_S_1503_out0 = v_S_9453_out0;
assign v_G1_4055_out0 = v_CARRY_4988_out0 || v_CARRY_4987_out0;
assign v_G1_4279_out0 = v_CARRY_5452_out0 || v_CARRY_5451_out0;
assign v_COUT_747_out0 = v_G1_4055_out0;
assign v_COUT_971_out0 = v_G1_4279_out0;
assign v__4553_out0 = { v__1829_out0,v_S_1279_out0 };
assign v__4568_out0 = { v__1844_out0,v_S_1503_out0 };
assign v_RM_3416_out0 = v_COUT_747_out0;
assign v_RM_3640_out0 = v_COUT_971_out0;
assign v_RM_11429_out0 = v_RM_3416_out0;
assign v_RM_11893_out0 = v_RM_3640_out0;
assign v_G1_7844_out0 = ((v_RD_5989_out0 && !v_RM_11429_out0) || (!v_RD_5989_out0) && v_RM_11429_out0);
assign v_G1_8308_out0 = ((v_RD_6453_out0 && !v_RM_11893_out0) || (!v_RD_6453_out0) && v_RM_11893_out0);
assign v_G2_12380_out0 = v_RD_5989_out0 && v_RM_11429_out0;
assign v_G2_12844_out0 = v_RD_6453_out0 && v_RM_11893_out0;
assign v_CARRY_4989_out0 = v_G2_12380_out0;
assign v_CARRY_5453_out0 = v_G2_12844_out0;
assign v_S_8990_out0 = v_G1_7844_out0;
assign v_S_9454_out0 = v_G1_8308_out0;
assign v_RM_11430_out0 = v_S_8990_out0;
assign v_RM_11894_out0 = v_S_9454_out0;
assign v_G1_7845_out0 = ((v_RD_5990_out0 && !v_RM_11430_out0) || (!v_RD_5990_out0) && v_RM_11430_out0);
assign v_G1_8309_out0 = ((v_RD_6454_out0 && !v_RM_11894_out0) || (!v_RD_6454_out0) && v_RM_11894_out0);
assign v_G2_12381_out0 = v_RD_5990_out0 && v_RM_11430_out0;
assign v_G2_12845_out0 = v_RD_6454_out0 && v_RM_11894_out0;
assign v_CARRY_4990_out0 = v_G2_12381_out0;
assign v_CARRY_5454_out0 = v_G2_12845_out0;
assign v_S_8991_out0 = v_G1_7845_out0;
assign v_S_9455_out0 = v_G1_8309_out0;
assign v_S_1280_out0 = v_S_8991_out0;
assign v_S_1504_out0 = v_S_9455_out0;
assign v_G1_4056_out0 = v_CARRY_4990_out0 || v_CARRY_4989_out0;
assign v_G1_4280_out0 = v_CARRY_5454_out0 || v_CARRY_5453_out0;
assign v_COUT_748_out0 = v_G1_4056_out0;
assign v_COUT_972_out0 = v_G1_4280_out0;
assign v__10655_out0 = { v__4553_out0,v_S_1280_out0 };
assign v__10670_out0 = { v__4568_out0,v_S_1504_out0 };
assign v__10950_out0 = { v__10655_out0,v_COUT_748_out0 };
assign v__10965_out0 = { v__10670_out0,v_COUT_972_out0 };
assign v_COUT_10920_out0 = v__10950_out0;
assign v_COUT_10935_out0 = v__10965_out0;
assign v_CIN_2355_out0 = v_COUT_10920_out0;
assign v_CIN_2370_out0 = v_COUT_10935_out0;
assign v__468_out0 = v_CIN_2355_out0[8:8];
assign v__483_out0 = v_CIN_2370_out0[8:8];
assign v__1773_out0 = v_CIN_2355_out0[6:6];
assign v__1788_out0 = v_CIN_2370_out0[6:6];
assign v__2155_out0 = v_CIN_2355_out0[3:3];
assign v__2170_out0 = v_CIN_2370_out0[3:3];
assign v__2195_out0 = v_CIN_2355_out0[15:15];
assign v__2209_out0 = v_CIN_2370_out0[15:15];
assign v__2502_out0 = v_CIN_2355_out0[0:0];
assign v__2517_out0 = v_CIN_2370_out0[0:0];
assign v__3051_out0 = v_CIN_2355_out0[9:9];
assign v__3066_out0 = v_CIN_2370_out0[9:9];
assign v__3085_out0 = v_CIN_2355_out0[2:2];
assign v__3100_out0 = v_CIN_2370_out0[2:2];
assign v__3139_out0 = v_CIN_2355_out0[7:7];
assign v__3154_out0 = v_CIN_2370_out0[7:7];
assign v__3823_out0 = v_CIN_2355_out0[1:1];
assign v__3838_out0 = v_CIN_2370_out0[1:1];
assign v__3861_out0 = v_CIN_2355_out0[10:10];
assign v__3876_out0 = v_CIN_2370_out0[10:10];
assign v__6800_out0 = v_CIN_2355_out0[11:11];
assign v__6815_out0 = v_CIN_2370_out0[11:11];
assign v__7644_out0 = v_CIN_2355_out0[12:12];
assign v__7659_out0 = v_CIN_2370_out0[12:12];
assign v__8699_out0 = v_CIN_2355_out0[13:13];
assign v__8714_out0 = v_CIN_2370_out0[13:13];
assign v__8769_out0 = v_CIN_2355_out0[14:14];
assign v__8784_out0 = v_CIN_2370_out0[14:14];
assign v__10719_out0 = v_CIN_2355_out0[5:5];
assign v__10734_out0 = v_CIN_2370_out0[5:5];
assign v__13448_out0 = v_CIN_2355_out0[4:4];
assign v__13463_out0 = v_CIN_2370_out0[4:4];
assign v_RM_3355_out0 = v__7644_out0;
assign v_RM_3356_out0 = v__8769_out0;
assign v_RM_3358_out0 = v__10719_out0;
assign v_RM_3359_out0 = v__13448_out0;
assign v_RM_3360_out0 = v__8699_out0;
assign v_RM_3361_out0 = v__3051_out0;
assign v_RM_3362_out0 = v__3861_out0;
assign v_RM_3363_out0 = v__3823_out0;
assign v_RM_3364_out0 = v__2155_out0;
assign v_RM_3365_out0 = v__1773_out0;
assign v_RM_3366_out0 = v__3139_out0;
assign v_RM_3367_out0 = v__6800_out0;
assign v_RM_3368_out0 = v__468_out0;
assign v_RM_3369_out0 = v__3085_out0;
assign v_RM_3579_out0 = v__7659_out0;
assign v_RM_3580_out0 = v__8784_out0;
assign v_RM_3582_out0 = v__10734_out0;
assign v_RM_3583_out0 = v__13463_out0;
assign v_RM_3584_out0 = v__8714_out0;
assign v_RM_3585_out0 = v__3066_out0;
assign v_RM_3586_out0 = v__3876_out0;
assign v_RM_3587_out0 = v__3838_out0;
assign v_RM_3588_out0 = v__2170_out0;
assign v_RM_3589_out0 = v__1788_out0;
assign v_RM_3590_out0 = v__3154_out0;
assign v_RM_3591_out0 = v__6815_out0;
assign v_RM_3592_out0 = v__483_out0;
assign v_RM_3593_out0 = v__3100_out0;
assign v_CIN_9810_out0 = v__2195_out0;
assign v_CIN_10034_out0 = v__2209_out0;
assign v_RM_11314_out0 = v__2502_out0;
assign v_RM_11778_out0 = v__2517_out0;
assign v_RD_5867_out0 = v_CIN_9810_out0;
assign v_RD_6331_out0 = v_CIN_10034_out0;
assign v_G1_7729_out0 = ((v_RD_5874_out0 && !v_RM_11314_out0) || (!v_RD_5874_out0) && v_RM_11314_out0);
assign v_G1_8193_out0 = ((v_RD_6338_out0 && !v_RM_11778_out0) || (!v_RD_6338_out0) && v_RM_11778_out0);
assign v_RM_11302_out0 = v_RM_3355_out0;
assign v_RM_11304_out0 = v_RM_3356_out0;
assign v_RM_11308_out0 = v_RM_3358_out0;
assign v_RM_11310_out0 = v_RM_3359_out0;
assign v_RM_11312_out0 = v_RM_3360_out0;
assign v_RM_11315_out0 = v_RM_3361_out0;
assign v_RM_11317_out0 = v_RM_3362_out0;
assign v_RM_11319_out0 = v_RM_3363_out0;
assign v_RM_11321_out0 = v_RM_3364_out0;
assign v_RM_11323_out0 = v_RM_3365_out0;
assign v_RM_11325_out0 = v_RM_3366_out0;
assign v_RM_11327_out0 = v_RM_3367_out0;
assign v_RM_11329_out0 = v_RM_3368_out0;
assign v_RM_11331_out0 = v_RM_3369_out0;
assign v_RM_11766_out0 = v_RM_3579_out0;
assign v_RM_11768_out0 = v_RM_3580_out0;
assign v_RM_11772_out0 = v_RM_3582_out0;
assign v_RM_11774_out0 = v_RM_3583_out0;
assign v_RM_11776_out0 = v_RM_3584_out0;
assign v_RM_11779_out0 = v_RM_3585_out0;
assign v_RM_11781_out0 = v_RM_3586_out0;
assign v_RM_11783_out0 = v_RM_3587_out0;
assign v_RM_11785_out0 = v_RM_3588_out0;
assign v_RM_11787_out0 = v_RM_3589_out0;
assign v_RM_11789_out0 = v_RM_3590_out0;
assign v_RM_11791_out0 = v_RM_3591_out0;
assign v_RM_11793_out0 = v_RM_3592_out0;
assign v_RM_11795_out0 = v_RM_3593_out0;
assign v_G2_12265_out0 = v_RD_5874_out0 && v_RM_11314_out0;
assign v_G2_12729_out0 = v_RD_6338_out0 && v_RM_11778_out0;
assign v_CARRY_4874_out0 = v_G2_12265_out0;
assign v_CARRY_5338_out0 = v_G2_12729_out0;
assign v_G1_7717_out0 = ((v_RD_5862_out0 && !v_RM_11302_out0) || (!v_RD_5862_out0) && v_RM_11302_out0);
assign v_G1_7719_out0 = ((v_RD_5864_out0 && !v_RM_11304_out0) || (!v_RD_5864_out0) && v_RM_11304_out0);
assign v_G1_7723_out0 = ((v_RD_5868_out0 && !v_RM_11308_out0) || (!v_RD_5868_out0) && v_RM_11308_out0);
assign v_G1_7725_out0 = ((v_RD_5870_out0 && !v_RM_11310_out0) || (!v_RD_5870_out0) && v_RM_11310_out0);
assign v_G1_7727_out0 = ((v_RD_5872_out0 && !v_RM_11312_out0) || (!v_RD_5872_out0) && v_RM_11312_out0);
assign v_G1_7730_out0 = ((v_RD_5875_out0 && !v_RM_11315_out0) || (!v_RD_5875_out0) && v_RM_11315_out0);
assign v_G1_7732_out0 = ((v_RD_5877_out0 && !v_RM_11317_out0) || (!v_RD_5877_out0) && v_RM_11317_out0);
assign v_G1_7734_out0 = ((v_RD_5879_out0 && !v_RM_11319_out0) || (!v_RD_5879_out0) && v_RM_11319_out0);
assign v_G1_7736_out0 = ((v_RD_5881_out0 && !v_RM_11321_out0) || (!v_RD_5881_out0) && v_RM_11321_out0);
assign v_G1_7738_out0 = ((v_RD_5883_out0 && !v_RM_11323_out0) || (!v_RD_5883_out0) && v_RM_11323_out0);
assign v_G1_7740_out0 = ((v_RD_5885_out0 && !v_RM_11325_out0) || (!v_RD_5885_out0) && v_RM_11325_out0);
assign v_G1_7742_out0 = ((v_RD_5887_out0 && !v_RM_11327_out0) || (!v_RD_5887_out0) && v_RM_11327_out0);
assign v_G1_7744_out0 = ((v_RD_5889_out0 && !v_RM_11329_out0) || (!v_RD_5889_out0) && v_RM_11329_out0);
assign v_G1_7746_out0 = ((v_RD_5891_out0 && !v_RM_11331_out0) || (!v_RD_5891_out0) && v_RM_11331_out0);
assign v_G1_8181_out0 = ((v_RD_6326_out0 && !v_RM_11766_out0) || (!v_RD_6326_out0) && v_RM_11766_out0);
assign v_G1_8183_out0 = ((v_RD_6328_out0 && !v_RM_11768_out0) || (!v_RD_6328_out0) && v_RM_11768_out0);
assign v_G1_8187_out0 = ((v_RD_6332_out0 && !v_RM_11772_out0) || (!v_RD_6332_out0) && v_RM_11772_out0);
assign v_G1_8189_out0 = ((v_RD_6334_out0 && !v_RM_11774_out0) || (!v_RD_6334_out0) && v_RM_11774_out0);
assign v_G1_8191_out0 = ((v_RD_6336_out0 && !v_RM_11776_out0) || (!v_RD_6336_out0) && v_RM_11776_out0);
assign v_G1_8194_out0 = ((v_RD_6339_out0 && !v_RM_11779_out0) || (!v_RD_6339_out0) && v_RM_11779_out0);
assign v_G1_8196_out0 = ((v_RD_6341_out0 && !v_RM_11781_out0) || (!v_RD_6341_out0) && v_RM_11781_out0);
assign v_G1_8198_out0 = ((v_RD_6343_out0 && !v_RM_11783_out0) || (!v_RD_6343_out0) && v_RM_11783_out0);
assign v_G1_8200_out0 = ((v_RD_6345_out0 && !v_RM_11785_out0) || (!v_RD_6345_out0) && v_RM_11785_out0);
assign v_G1_8202_out0 = ((v_RD_6347_out0 && !v_RM_11787_out0) || (!v_RD_6347_out0) && v_RM_11787_out0);
assign v_G1_8204_out0 = ((v_RD_6349_out0 && !v_RM_11789_out0) || (!v_RD_6349_out0) && v_RM_11789_out0);
assign v_G1_8206_out0 = ((v_RD_6351_out0 && !v_RM_11791_out0) || (!v_RD_6351_out0) && v_RM_11791_out0);
assign v_G1_8208_out0 = ((v_RD_6353_out0 && !v_RM_11793_out0) || (!v_RD_6353_out0) && v_RM_11793_out0);
assign v_G1_8210_out0 = ((v_RD_6355_out0 && !v_RM_11795_out0) || (!v_RD_6355_out0) && v_RM_11795_out0);
assign v_S_8875_out0 = v_G1_7729_out0;
assign v_S_9339_out0 = v_G1_8193_out0;
assign v_G2_12253_out0 = v_RD_5862_out0 && v_RM_11302_out0;
assign v_G2_12255_out0 = v_RD_5864_out0 && v_RM_11304_out0;
assign v_G2_12259_out0 = v_RD_5868_out0 && v_RM_11308_out0;
assign v_G2_12261_out0 = v_RD_5870_out0 && v_RM_11310_out0;
assign v_G2_12263_out0 = v_RD_5872_out0 && v_RM_11312_out0;
assign v_G2_12266_out0 = v_RD_5875_out0 && v_RM_11315_out0;
assign v_G2_12268_out0 = v_RD_5877_out0 && v_RM_11317_out0;
assign v_G2_12270_out0 = v_RD_5879_out0 && v_RM_11319_out0;
assign v_G2_12272_out0 = v_RD_5881_out0 && v_RM_11321_out0;
assign v_G2_12274_out0 = v_RD_5883_out0 && v_RM_11323_out0;
assign v_G2_12276_out0 = v_RD_5885_out0 && v_RM_11325_out0;
assign v_G2_12278_out0 = v_RD_5887_out0 && v_RM_11327_out0;
assign v_G2_12280_out0 = v_RD_5889_out0 && v_RM_11329_out0;
assign v_G2_12282_out0 = v_RD_5891_out0 && v_RM_11331_out0;
assign v_G2_12717_out0 = v_RD_6326_out0 && v_RM_11766_out0;
assign v_G2_12719_out0 = v_RD_6328_out0 && v_RM_11768_out0;
assign v_G2_12723_out0 = v_RD_6332_out0 && v_RM_11772_out0;
assign v_G2_12725_out0 = v_RD_6334_out0 && v_RM_11774_out0;
assign v_G2_12727_out0 = v_RD_6336_out0 && v_RM_11776_out0;
assign v_G2_12730_out0 = v_RD_6339_out0 && v_RM_11779_out0;
assign v_G2_12732_out0 = v_RD_6341_out0 && v_RM_11781_out0;
assign v_G2_12734_out0 = v_RD_6343_out0 && v_RM_11783_out0;
assign v_G2_12736_out0 = v_RD_6345_out0 && v_RM_11785_out0;
assign v_G2_12738_out0 = v_RD_6347_out0 && v_RM_11787_out0;
assign v_G2_12740_out0 = v_RD_6349_out0 && v_RM_11789_out0;
assign v_G2_12742_out0 = v_RD_6351_out0 && v_RM_11791_out0;
assign v_G2_12744_out0 = v_RD_6353_out0 && v_RM_11793_out0;
assign v_G2_12746_out0 = v_RD_6355_out0 && v_RM_11795_out0;
assign v_S_4665_out0 = v_S_8875_out0;
assign v_S_4680_out0 = v_S_9339_out0;
assign v_CARRY_4862_out0 = v_G2_12253_out0;
assign v_CARRY_4864_out0 = v_G2_12255_out0;
assign v_CARRY_4868_out0 = v_G2_12259_out0;
assign v_CARRY_4870_out0 = v_G2_12261_out0;
assign v_CARRY_4872_out0 = v_G2_12263_out0;
assign v_CARRY_4875_out0 = v_G2_12266_out0;
assign v_CARRY_4877_out0 = v_G2_12268_out0;
assign v_CARRY_4879_out0 = v_G2_12270_out0;
assign v_CARRY_4881_out0 = v_G2_12272_out0;
assign v_CARRY_4883_out0 = v_G2_12274_out0;
assign v_CARRY_4885_out0 = v_G2_12276_out0;
assign v_CARRY_4887_out0 = v_G2_12278_out0;
assign v_CARRY_4889_out0 = v_G2_12280_out0;
assign v_CARRY_4891_out0 = v_G2_12282_out0;
assign v_CARRY_5326_out0 = v_G2_12717_out0;
assign v_CARRY_5328_out0 = v_G2_12719_out0;
assign v_CARRY_5332_out0 = v_G2_12723_out0;
assign v_CARRY_5334_out0 = v_G2_12725_out0;
assign v_CARRY_5336_out0 = v_G2_12727_out0;
assign v_CARRY_5339_out0 = v_G2_12730_out0;
assign v_CARRY_5341_out0 = v_G2_12732_out0;
assign v_CARRY_5343_out0 = v_G2_12734_out0;
assign v_CARRY_5345_out0 = v_G2_12736_out0;
assign v_CARRY_5347_out0 = v_G2_12738_out0;
assign v_CARRY_5349_out0 = v_G2_12740_out0;
assign v_CARRY_5351_out0 = v_G2_12742_out0;
assign v_CARRY_5353_out0 = v_G2_12744_out0;
assign v_CARRY_5355_out0 = v_G2_12746_out0;
assign v_S_8863_out0 = v_G1_7717_out0;
assign v_S_8865_out0 = v_G1_7719_out0;
assign v_S_8869_out0 = v_G1_7723_out0;
assign v_S_8871_out0 = v_G1_7725_out0;
assign v_S_8873_out0 = v_G1_7727_out0;
assign v_S_8876_out0 = v_G1_7730_out0;
assign v_S_8878_out0 = v_G1_7732_out0;
assign v_S_8880_out0 = v_G1_7734_out0;
assign v_S_8882_out0 = v_G1_7736_out0;
assign v_S_8884_out0 = v_G1_7738_out0;
assign v_S_8886_out0 = v_G1_7740_out0;
assign v_S_8888_out0 = v_G1_7742_out0;
assign v_S_8890_out0 = v_G1_7744_out0;
assign v_S_8892_out0 = v_G1_7746_out0;
assign v_S_9327_out0 = v_G1_8181_out0;
assign v_S_9329_out0 = v_G1_8183_out0;
assign v_S_9333_out0 = v_G1_8187_out0;
assign v_S_9335_out0 = v_G1_8189_out0;
assign v_S_9337_out0 = v_G1_8191_out0;
assign v_S_9340_out0 = v_G1_8194_out0;
assign v_S_9342_out0 = v_G1_8196_out0;
assign v_S_9344_out0 = v_G1_8198_out0;
assign v_S_9346_out0 = v_G1_8200_out0;
assign v_S_9348_out0 = v_G1_8202_out0;
assign v_S_9350_out0 = v_G1_8204_out0;
assign v_S_9352_out0 = v_G1_8206_out0;
assign v_S_9354_out0 = v_G1_8208_out0;
assign v_S_9356_out0 = v_G1_8210_out0;
assign v_CIN_9816_out0 = v_CARRY_4874_out0;
assign v_CIN_10040_out0 = v_CARRY_5338_out0;
assign v__2392_out0 = { v__4529_out0,v_S_4665_out0 };
assign v__2393_out0 = { v__4530_out0,v_S_4680_out0 };
assign v_RD_5880_out0 = v_CIN_9816_out0;
assign v_RD_6344_out0 = v_CIN_10040_out0;
assign v_RM_11303_out0 = v_S_8863_out0;
assign v_RM_11305_out0 = v_S_8865_out0;
assign v_RM_11309_out0 = v_S_8869_out0;
assign v_RM_11311_out0 = v_S_8871_out0;
assign v_RM_11313_out0 = v_S_8873_out0;
assign v_RM_11316_out0 = v_S_8876_out0;
assign v_RM_11318_out0 = v_S_8878_out0;
assign v_RM_11320_out0 = v_S_8880_out0;
assign v_RM_11322_out0 = v_S_8882_out0;
assign v_RM_11324_out0 = v_S_8884_out0;
assign v_RM_11326_out0 = v_S_8886_out0;
assign v_RM_11328_out0 = v_S_8888_out0;
assign v_RM_11330_out0 = v_S_8890_out0;
assign v_RM_11332_out0 = v_S_8892_out0;
assign v_RM_11767_out0 = v_S_9327_out0;
assign v_RM_11769_out0 = v_S_9329_out0;
assign v_RM_11773_out0 = v_S_9333_out0;
assign v_RM_11775_out0 = v_S_9335_out0;
assign v_RM_11777_out0 = v_S_9337_out0;
assign v_RM_11780_out0 = v_S_9340_out0;
assign v_RM_11782_out0 = v_S_9342_out0;
assign v_RM_11784_out0 = v_S_9344_out0;
assign v_RM_11786_out0 = v_S_9346_out0;
assign v_RM_11788_out0 = v_S_9348_out0;
assign v_RM_11790_out0 = v_S_9350_out0;
assign v_RM_11792_out0 = v_S_9352_out0;
assign v_RM_11794_out0 = v_S_9354_out0;
assign v_RM_11796_out0 = v_S_9356_out0;
assign v_G1_7735_out0 = ((v_RD_5880_out0 && !v_RM_11320_out0) || (!v_RD_5880_out0) && v_RM_11320_out0);
assign v_G1_8199_out0 = ((v_RD_6344_out0 && !v_RM_11784_out0) || (!v_RD_6344_out0) && v_RM_11784_out0);
assign v_G2_12271_out0 = v_RD_5880_out0 && v_RM_11320_out0;
assign v_G2_12735_out0 = v_RD_6344_out0 && v_RM_11784_out0;
assign v_CARRY_4880_out0 = v_G2_12271_out0;
assign v_CARRY_5344_out0 = v_G2_12735_out0;
assign v_S_8881_out0 = v_G1_7735_out0;
assign v_S_9345_out0 = v_G1_8199_out0;
assign v_S_1227_out0 = v_S_8881_out0;
assign v_S_1451_out0 = v_S_9345_out0;
assign v_G1_4003_out0 = v_CARRY_4880_out0 || v_CARRY_4879_out0;
assign v_G1_4227_out0 = v_CARRY_5344_out0 || v_CARRY_5343_out0;
assign v_COUT_695_out0 = v_G1_4003_out0;
assign v_COUT_919_out0 = v_G1_4227_out0;
assign v_CIN_9822_out0 = v_COUT_695_out0;
assign v_CIN_10046_out0 = v_COUT_919_out0;
assign v_RD_5892_out0 = v_CIN_9822_out0;
assign v_RD_6356_out0 = v_CIN_10046_out0;
assign v_G1_7747_out0 = ((v_RD_5892_out0 && !v_RM_11332_out0) || (!v_RD_5892_out0) && v_RM_11332_out0);
assign v_G1_8211_out0 = ((v_RD_6356_out0 && !v_RM_11796_out0) || (!v_RD_6356_out0) && v_RM_11796_out0);
assign v_G2_12283_out0 = v_RD_5892_out0 && v_RM_11332_out0;
assign v_G2_12747_out0 = v_RD_6356_out0 && v_RM_11796_out0;
assign v_CARRY_4892_out0 = v_G2_12283_out0;
assign v_CARRY_5356_out0 = v_G2_12747_out0;
assign v_S_8893_out0 = v_G1_7747_out0;
assign v_S_9357_out0 = v_G1_8211_out0;
assign v_S_1233_out0 = v_S_8893_out0;
assign v_S_1457_out0 = v_S_9357_out0;
assign v_G1_4009_out0 = v_CARRY_4892_out0 || v_CARRY_4891_out0;
assign v_G1_4233_out0 = v_CARRY_5356_out0 || v_CARRY_5355_out0;
assign v_COUT_701_out0 = v_G1_4009_out0;
assign v_COUT_925_out0 = v_G1_4233_out0;
assign v__4782_out0 = { v_S_1227_out0,v_S_1233_out0 };
assign v__4797_out0 = { v_S_1451_out0,v_S_1457_out0 };
assign v_CIN_9817_out0 = v_COUT_701_out0;
assign v_CIN_10041_out0 = v_COUT_925_out0;
assign v_RD_5882_out0 = v_CIN_9817_out0;
assign v_RD_6346_out0 = v_CIN_10041_out0;
assign v_G1_7737_out0 = ((v_RD_5882_out0 && !v_RM_11322_out0) || (!v_RD_5882_out0) && v_RM_11322_out0);
assign v_G1_8201_out0 = ((v_RD_6346_out0 && !v_RM_11786_out0) || (!v_RD_6346_out0) && v_RM_11786_out0);
assign v_G2_12273_out0 = v_RD_5882_out0 && v_RM_11322_out0;
assign v_G2_12737_out0 = v_RD_6346_out0 && v_RM_11786_out0;
assign v_CARRY_4882_out0 = v_G2_12273_out0;
assign v_CARRY_5346_out0 = v_G2_12737_out0;
assign v_S_8883_out0 = v_G1_7737_out0;
assign v_S_9347_out0 = v_G1_8201_out0;
assign v_S_1228_out0 = v_S_8883_out0;
assign v_S_1452_out0 = v_S_9347_out0;
assign v_G1_4004_out0 = v_CARRY_4882_out0 || v_CARRY_4881_out0;
assign v_G1_4228_out0 = v_CARRY_5346_out0 || v_CARRY_5345_out0;
assign v_COUT_696_out0 = v_G1_4004_out0;
assign v_COUT_920_out0 = v_G1_4228_out0;
assign v__2552_out0 = { v__4782_out0,v_S_1228_out0 };
assign v__2567_out0 = { v__4797_out0,v_S_1452_out0 };
assign v_CIN_9812_out0 = v_COUT_696_out0;
assign v_CIN_10036_out0 = v_COUT_920_out0;
assign v_RD_5871_out0 = v_CIN_9812_out0;
assign v_RD_6335_out0 = v_CIN_10036_out0;
assign v_G1_7726_out0 = ((v_RD_5871_out0 && !v_RM_11311_out0) || (!v_RD_5871_out0) && v_RM_11311_out0);
assign v_G1_8190_out0 = ((v_RD_6335_out0 && !v_RM_11775_out0) || (!v_RD_6335_out0) && v_RM_11775_out0);
assign v_G2_12262_out0 = v_RD_5871_out0 && v_RM_11311_out0;
assign v_G2_12726_out0 = v_RD_6335_out0 && v_RM_11775_out0;
assign v_CARRY_4871_out0 = v_G2_12262_out0;
assign v_CARRY_5335_out0 = v_G2_12726_out0;
assign v_S_8872_out0 = v_G1_7726_out0;
assign v_S_9336_out0 = v_G1_8190_out0;
assign v_S_1223_out0 = v_S_8872_out0;
assign v_S_1447_out0 = v_S_9336_out0;
assign v_G1_3999_out0 = v_CARRY_4871_out0 || v_CARRY_4870_out0;
assign v_G1_4223_out0 = v_CARRY_5335_out0 || v_CARRY_5334_out0;
assign v_COUT_691_out0 = v_G1_3999_out0;
assign v_COUT_915_out0 = v_G1_4223_out0;
assign v__7032_out0 = { v__2552_out0,v_S_1223_out0 };
assign v__7047_out0 = { v__2567_out0,v_S_1447_out0 };
assign v_CIN_9811_out0 = v_COUT_691_out0;
assign v_CIN_10035_out0 = v_COUT_915_out0;
assign v_RD_5869_out0 = v_CIN_9811_out0;
assign v_RD_6333_out0 = v_CIN_10035_out0;
assign v_G1_7724_out0 = ((v_RD_5869_out0 && !v_RM_11309_out0) || (!v_RD_5869_out0) && v_RM_11309_out0);
assign v_G1_8188_out0 = ((v_RD_6333_out0 && !v_RM_11773_out0) || (!v_RD_6333_out0) && v_RM_11773_out0);
assign v_G2_12260_out0 = v_RD_5869_out0 && v_RM_11309_out0;
assign v_G2_12724_out0 = v_RD_6333_out0 && v_RM_11773_out0;
assign v_CARRY_4869_out0 = v_G2_12260_out0;
assign v_CARRY_5333_out0 = v_G2_12724_out0;
assign v_S_8870_out0 = v_G1_7724_out0;
assign v_S_9334_out0 = v_G1_8188_out0;
assign v_S_1222_out0 = v_S_8870_out0;
assign v_S_1446_out0 = v_S_9334_out0;
assign v_G1_3998_out0 = v_CARRY_4869_out0 || v_CARRY_4868_out0;
assign v_G1_4222_out0 = v_CARRY_5333_out0 || v_CARRY_5332_out0;
assign v_COUT_690_out0 = v_G1_3998_out0;
assign v_COUT_914_out0 = v_G1_4222_out0;
assign v__13518_out0 = { v__7032_out0,v_S_1222_out0 };
assign v__13533_out0 = { v__7047_out0,v_S_1446_out0 };
assign v_CIN_9818_out0 = v_COUT_690_out0;
assign v_CIN_10042_out0 = v_COUT_914_out0;
assign v_RD_5884_out0 = v_CIN_9818_out0;
assign v_RD_6348_out0 = v_CIN_10042_out0;
assign v_G1_7739_out0 = ((v_RD_5884_out0 && !v_RM_11324_out0) || (!v_RD_5884_out0) && v_RM_11324_out0);
assign v_G1_8203_out0 = ((v_RD_6348_out0 && !v_RM_11788_out0) || (!v_RD_6348_out0) && v_RM_11788_out0);
assign v_G2_12275_out0 = v_RD_5884_out0 && v_RM_11324_out0;
assign v_G2_12739_out0 = v_RD_6348_out0 && v_RM_11788_out0;
assign v_CARRY_4884_out0 = v_G2_12275_out0;
assign v_CARRY_5348_out0 = v_G2_12739_out0;
assign v_S_8885_out0 = v_G1_7739_out0;
assign v_S_9349_out0 = v_G1_8203_out0;
assign v_S_1229_out0 = v_S_8885_out0;
assign v_S_1453_out0 = v_S_9349_out0;
assign v_G1_4005_out0 = v_CARRY_4884_out0 || v_CARRY_4883_out0;
assign v_G1_4229_out0 = v_CARRY_5348_out0 || v_CARRY_5347_out0;
assign v_COUT_697_out0 = v_G1_4005_out0;
assign v_COUT_921_out0 = v_G1_4229_out0;
assign v__3311_out0 = { v__13518_out0,v_S_1229_out0 };
assign v__3326_out0 = { v__13533_out0,v_S_1453_out0 };
assign v_CIN_9819_out0 = v_COUT_697_out0;
assign v_CIN_10043_out0 = v_COUT_921_out0;
assign v_RD_5886_out0 = v_CIN_9819_out0;
assign v_RD_6350_out0 = v_CIN_10043_out0;
assign v_G1_7741_out0 = ((v_RD_5886_out0 && !v_RM_11326_out0) || (!v_RD_5886_out0) && v_RM_11326_out0);
assign v_G1_8205_out0 = ((v_RD_6350_out0 && !v_RM_11790_out0) || (!v_RD_6350_out0) && v_RM_11790_out0);
assign v_G2_12277_out0 = v_RD_5886_out0 && v_RM_11326_out0;
assign v_G2_12741_out0 = v_RD_6350_out0 && v_RM_11790_out0;
assign v_CARRY_4886_out0 = v_G2_12277_out0;
assign v_CARRY_5350_out0 = v_G2_12741_out0;
assign v_S_8887_out0 = v_G1_7741_out0;
assign v_S_9351_out0 = v_G1_8205_out0;
assign v_S_1230_out0 = v_S_8887_out0;
assign v_S_1454_out0 = v_S_9351_out0;
assign v_G1_4006_out0 = v_CARRY_4886_out0 || v_CARRY_4885_out0;
assign v_G1_4230_out0 = v_CARRY_5350_out0 || v_CARRY_5349_out0;
assign v_COUT_698_out0 = v_G1_4006_out0;
assign v_COUT_922_out0 = v_G1_4230_out0;
assign v__7147_out0 = { v__3311_out0,v_S_1230_out0 };
assign v__7162_out0 = { v__3326_out0,v_S_1454_out0 };
assign v_CIN_9821_out0 = v_COUT_698_out0;
assign v_CIN_10045_out0 = v_COUT_922_out0;
assign v_RD_5890_out0 = v_CIN_9821_out0;
assign v_RD_6354_out0 = v_CIN_10045_out0;
assign v_G1_7745_out0 = ((v_RD_5890_out0 && !v_RM_11330_out0) || (!v_RD_5890_out0) && v_RM_11330_out0);
assign v_G1_8209_out0 = ((v_RD_6354_out0 && !v_RM_11794_out0) || (!v_RD_6354_out0) && v_RM_11794_out0);
assign v_G2_12281_out0 = v_RD_5890_out0 && v_RM_11330_out0;
assign v_G2_12745_out0 = v_RD_6354_out0 && v_RM_11794_out0;
assign v_CARRY_4890_out0 = v_G2_12281_out0;
assign v_CARRY_5354_out0 = v_G2_12745_out0;
assign v_S_8891_out0 = v_G1_7745_out0;
assign v_S_9355_out0 = v_G1_8209_out0;
assign v_S_1232_out0 = v_S_8891_out0;
assign v_S_1456_out0 = v_S_9355_out0;
assign v_G1_4008_out0 = v_CARRY_4890_out0 || v_CARRY_4889_out0;
assign v_G1_4232_out0 = v_CARRY_5354_out0 || v_CARRY_5353_out0;
assign v_COUT_700_out0 = v_G1_4008_out0;
assign v_COUT_924_out0 = v_G1_4232_out0;
assign v__4749_out0 = { v__7147_out0,v_S_1232_out0 };
assign v__4764_out0 = { v__7162_out0,v_S_1456_out0 };
assign v_CIN_9814_out0 = v_COUT_700_out0;
assign v_CIN_10038_out0 = v_COUT_924_out0;
assign v_RD_5876_out0 = v_CIN_9814_out0;
assign v_RD_6340_out0 = v_CIN_10038_out0;
assign v_G1_7731_out0 = ((v_RD_5876_out0 && !v_RM_11316_out0) || (!v_RD_5876_out0) && v_RM_11316_out0);
assign v_G1_8195_out0 = ((v_RD_6340_out0 && !v_RM_11780_out0) || (!v_RD_6340_out0) && v_RM_11780_out0);
assign v_G2_12267_out0 = v_RD_5876_out0 && v_RM_11316_out0;
assign v_G2_12731_out0 = v_RD_6340_out0 && v_RM_11780_out0;
assign v_CARRY_4876_out0 = v_G2_12267_out0;
assign v_CARRY_5340_out0 = v_G2_12731_out0;
assign v_S_8877_out0 = v_G1_7731_out0;
assign v_S_9341_out0 = v_G1_8195_out0;
assign v_S_1225_out0 = v_S_8877_out0;
assign v_S_1449_out0 = v_S_9341_out0;
assign v_G1_4001_out0 = v_CARRY_4876_out0 || v_CARRY_4875_out0;
assign v_G1_4225_out0 = v_CARRY_5340_out0 || v_CARRY_5339_out0;
assign v_COUT_693_out0 = v_G1_4001_out0;
assign v_COUT_917_out0 = v_G1_4225_out0;
assign v__6926_out0 = { v__4749_out0,v_S_1225_out0 };
assign v__6941_out0 = { v__4764_out0,v_S_1449_out0 };
assign v_CIN_9815_out0 = v_COUT_693_out0;
assign v_CIN_10039_out0 = v_COUT_917_out0;
assign v_RD_5878_out0 = v_CIN_9815_out0;
assign v_RD_6342_out0 = v_CIN_10039_out0;
assign v_G1_7733_out0 = ((v_RD_5878_out0 && !v_RM_11318_out0) || (!v_RD_5878_out0) && v_RM_11318_out0);
assign v_G1_8197_out0 = ((v_RD_6342_out0 && !v_RM_11782_out0) || (!v_RD_6342_out0) && v_RM_11782_out0);
assign v_G2_12269_out0 = v_RD_5878_out0 && v_RM_11318_out0;
assign v_G2_12733_out0 = v_RD_6342_out0 && v_RM_11782_out0;
assign v_CARRY_4878_out0 = v_G2_12269_out0;
assign v_CARRY_5342_out0 = v_G2_12733_out0;
assign v_S_8879_out0 = v_G1_7733_out0;
assign v_S_9343_out0 = v_G1_8197_out0;
assign v_S_1226_out0 = v_S_8879_out0;
assign v_S_1450_out0 = v_S_9343_out0;
assign v_G1_4002_out0 = v_CARRY_4878_out0 || v_CARRY_4877_out0;
assign v_G1_4226_out0 = v_CARRY_5342_out0 || v_CARRY_5341_out0;
assign v_COUT_694_out0 = v_G1_4002_out0;
assign v_COUT_918_out0 = v_G1_4226_out0;
assign v__5802_out0 = { v__6926_out0,v_S_1226_out0 };
assign v__5817_out0 = { v__6941_out0,v_S_1450_out0 };
assign v_CIN_9820_out0 = v_COUT_694_out0;
assign v_CIN_10044_out0 = v_COUT_918_out0;
assign v_RD_5888_out0 = v_CIN_9820_out0;
assign v_RD_6352_out0 = v_CIN_10044_out0;
assign v_G1_7743_out0 = ((v_RD_5888_out0 && !v_RM_11328_out0) || (!v_RD_5888_out0) && v_RM_11328_out0);
assign v_G1_8207_out0 = ((v_RD_6352_out0 && !v_RM_11792_out0) || (!v_RD_6352_out0) && v_RM_11792_out0);
assign v_G2_12279_out0 = v_RD_5888_out0 && v_RM_11328_out0;
assign v_G2_12743_out0 = v_RD_6352_out0 && v_RM_11792_out0;
assign v_CARRY_4888_out0 = v_G2_12279_out0;
assign v_CARRY_5352_out0 = v_G2_12743_out0;
assign v_S_8889_out0 = v_G1_7743_out0;
assign v_S_9353_out0 = v_G1_8207_out0;
assign v_S_1231_out0 = v_S_8889_out0;
assign v_S_1455_out0 = v_S_9353_out0;
assign v_G1_4007_out0 = v_CARRY_4888_out0 || v_CARRY_4887_out0;
assign v_G1_4231_out0 = v_CARRY_5352_out0 || v_CARRY_5351_out0;
assign v_COUT_699_out0 = v_G1_4007_out0;
assign v_COUT_923_out0 = v_G1_4231_out0;
assign v__2026_out0 = { v__5802_out0,v_S_1231_out0 };
assign v__2041_out0 = { v__5817_out0,v_S_1455_out0 };
assign v_CIN_9808_out0 = v_COUT_699_out0;
assign v_CIN_10032_out0 = v_COUT_923_out0;
assign v_RD_5863_out0 = v_CIN_9808_out0;
assign v_RD_6327_out0 = v_CIN_10032_out0;
assign v_G1_7718_out0 = ((v_RD_5863_out0 && !v_RM_11303_out0) || (!v_RD_5863_out0) && v_RM_11303_out0);
assign v_G1_8182_out0 = ((v_RD_6327_out0 && !v_RM_11767_out0) || (!v_RD_6327_out0) && v_RM_11767_out0);
assign v_G2_12254_out0 = v_RD_5863_out0 && v_RM_11303_out0;
assign v_G2_12718_out0 = v_RD_6327_out0 && v_RM_11767_out0;
assign v_CARRY_4863_out0 = v_G2_12254_out0;
assign v_CARRY_5327_out0 = v_G2_12718_out0;
assign v_S_8864_out0 = v_G1_7718_out0;
assign v_S_9328_out0 = v_G1_8182_out0;
assign v_S_1219_out0 = v_S_8864_out0;
assign v_S_1443_out0 = v_S_9328_out0;
assign v_G1_3995_out0 = v_CARRY_4863_out0 || v_CARRY_4862_out0;
assign v_G1_4219_out0 = v_CARRY_5327_out0 || v_CARRY_5326_out0;
assign v_COUT_687_out0 = v_G1_3995_out0;
assign v_COUT_911_out0 = v_G1_4219_out0;
assign v__2793_out0 = { v__2026_out0,v_S_1219_out0 };
assign v__2808_out0 = { v__2041_out0,v_S_1443_out0 };
assign v_CIN_9813_out0 = v_COUT_687_out0;
assign v_CIN_10037_out0 = v_COUT_911_out0;
assign v_RD_5873_out0 = v_CIN_9813_out0;
assign v_RD_6337_out0 = v_CIN_10037_out0;
assign v_G1_7728_out0 = ((v_RD_5873_out0 && !v_RM_11313_out0) || (!v_RD_5873_out0) && v_RM_11313_out0);
assign v_G1_8192_out0 = ((v_RD_6337_out0 && !v_RM_11777_out0) || (!v_RD_6337_out0) && v_RM_11777_out0);
assign v_G2_12264_out0 = v_RD_5873_out0 && v_RM_11313_out0;
assign v_G2_12728_out0 = v_RD_6337_out0 && v_RM_11777_out0;
assign v_CARRY_4873_out0 = v_G2_12264_out0;
assign v_CARRY_5337_out0 = v_G2_12728_out0;
assign v_S_8874_out0 = v_G1_7728_out0;
assign v_S_9338_out0 = v_G1_8192_out0;
assign v_S_1224_out0 = v_S_8874_out0;
assign v_S_1448_out0 = v_S_9338_out0;
assign v_G1_4000_out0 = v_CARRY_4873_out0 || v_CARRY_4872_out0;
assign v_G1_4224_out0 = v_CARRY_5337_out0 || v_CARRY_5336_out0;
assign v_COUT_692_out0 = v_G1_4000_out0;
assign v_COUT_916_out0 = v_G1_4224_out0;
assign v__1825_out0 = { v__2793_out0,v_S_1224_out0 };
assign v__1840_out0 = { v__2808_out0,v_S_1448_out0 };
assign v_CIN_9809_out0 = v_COUT_692_out0;
assign v_CIN_10033_out0 = v_COUT_916_out0;
assign v_RD_5865_out0 = v_CIN_9809_out0;
assign v_RD_6329_out0 = v_CIN_10033_out0;
assign v_G1_7720_out0 = ((v_RD_5865_out0 && !v_RM_11305_out0) || (!v_RD_5865_out0) && v_RM_11305_out0);
assign v_G1_8184_out0 = ((v_RD_6329_out0 && !v_RM_11769_out0) || (!v_RD_6329_out0) && v_RM_11769_out0);
assign v_G2_12256_out0 = v_RD_5865_out0 && v_RM_11305_out0;
assign v_G2_12720_out0 = v_RD_6329_out0 && v_RM_11769_out0;
assign v_CARRY_4865_out0 = v_G2_12256_out0;
assign v_CARRY_5329_out0 = v_G2_12720_out0;
assign v_S_8866_out0 = v_G1_7720_out0;
assign v_S_9330_out0 = v_G1_8184_out0;
assign v_S_1220_out0 = v_S_8866_out0;
assign v_S_1444_out0 = v_S_9330_out0;
assign v_G1_3996_out0 = v_CARRY_4865_out0 || v_CARRY_4864_out0;
assign v_G1_4220_out0 = v_CARRY_5329_out0 || v_CARRY_5328_out0;
assign v_COUT_688_out0 = v_G1_3996_out0;
assign v_COUT_912_out0 = v_G1_4220_out0;
assign v__4549_out0 = { v__1825_out0,v_S_1220_out0 };
assign v__4564_out0 = { v__1840_out0,v_S_1444_out0 };
assign v_RM_3357_out0 = v_COUT_688_out0;
assign v_RM_3581_out0 = v_COUT_912_out0;
assign v_RM_11306_out0 = v_RM_3357_out0;
assign v_RM_11770_out0 = v_RM_3581_out0;
assign v_G1_7721_out0 = ((v_RD_5866_out0 && !v_RM_11306_out0) || (!v_RD_5866_out0) && v_RM_11306_out0);
assign v_G1_8185_out0 = ((v_RD_6330_out0 && !v_RM_11770_out0) || (!v_RD_6330_out0) && v_RM_11770_out0);
assign v_G2_12257_out0 = v_RD_5866_out0 && v_RM_11306_out0;
assign v_G2_12721_out0 = v_RD_6330_out0 && v_RM_11770_out0;
assign v_CARRY_4866_out0 = v_G2_12257_out0;
assign v_CARRY_5330_out0 = v_G2_12721_out0;
assign v_S_8867_out0 = v_G1_7721_out0;
assign v_S_9331_out0 = v_G1_8185_out0;
assign v_RM_11307_out0 = v_S_8867_out0;
assign v_RM_11771_out0 = v_S_9331_out0;
assign v_G1_7722_out0 = ((v_RD_5867_out0 && !v_RM_11307_out0) || (!v_RD_5867_out0) && v_RM_11307_out0);
assign v_G1_8186_out0 = ((v_RD_6331_out0 && !v_RM_11771_out0) || (!v_RD_6331_out0) && v_RM_11771_out0);
assign v_G2_12258_out0 = v_RD_5867_out0 && v_RM_11307_out0;
assign v_G2_12722_out0 = v_RD_6331_out0 && v_RM_11771_out0;
assign v_CARRY_4867_out0 = v_G2_12258_out0;
assign v_CARRY_5331_out0 = v_G2_12722_out0;
assign v_S_8868_out0 = v_G1_7722_out0;
assign v_S_9332_out0 = v_G1_8186_out0;
assign v_S_1221_out0 = v_S_8868_out0;
assign v_S_1445_out0 = v_S_9332_out0;
assign v_G1_3997_out0 = v_CARRY_4867_out0 || v_CARRY_4866_out0;
assign v_G1_4221_out0 = v_CARRY_5331_out0 || v_CARRY_5330_out0;
assign v_COUT_689_out0 = v_G1_3997_out0;
assign v_COUT_913_out0 = v_G1_4221_out0;
assign v__10651_out0 = { v__4549_out0,v_S_1221_out0 };
assign v__10666_out0 = { v__4564_out0,v_S_1445_out0 };
assign v__10946_out0 = { v__10651_out0,v_COUT_689_out0 };
assign v__10961_out0 = { v__10666_out0,v_COUT_913_out0 };
assign v_COUT_10916_out0 = v__10946_out0;
assign v_COUT_10931_out0 = v__10961_out0;
assign v_CIN_2365_out0 = v_COUT_10916_out0;
assign v_CIN_2380_out0 = v_COUT_10931_out0;
assign v__478_out0 = v_CIN_2365_out0[8:8];
assign v__493_out0 = v_CIN_2380_out0[8:8];
assign v__1783_out0 = v_CIN_2365_out0[6:6];
assign v__1798_out0 = v_CIN_2380_out0[6:6];
assign v__2165_out0 = v_CIN_2365_out0[3:3];
assign v__2180_out0 = v_CIN_2380_out0[3:3];
assign v__2204_out0 = v_CIN_2365_out0[15:15];
assign v__2218_out0 = v_CIN_2380_out0[15:15];
assign v__2512_out0 = v_CIN_2365_out0[0:0];
assign v__2527_out0 = v_CIN_2380_out0[0:0];
assign v__3061_out0 = v_CIN_2365_out0[9:9];
assign v__3076_out0 = v_CIN_2380_out0[9:9];
assign v__3095_out0 = v_CIN_2365_out0[2:2];
assign v__3110_out0 = v_CIN_2380_out0[2:2];
assign v__3149_out0 = v_CIN_2365_out0[7:7];
assign v__3164_out0 = v_CIN_2380_out0[7:7];
assign v__3833_out0 = v_CIN_2365_out0[1:1];
assign v__3848_out0 = v_CIN_2380_out0[1:1];
assign v__3871_out0 = v_CIN_2365_out0[10:10];
assign v__3886_out0 = v_CIN_2380_out0[10:10];
assign v__6810_out0 = v_CIN_2365_out0[11:11];
assign v__6825_out0 = v_CIN_2380_out0[11:11];
assign v__7654_out0 = v_CIN_2365_out0[12:12];
assign v__7669_out0 = v_CIN_2380_out0[12:12];
assign v__8709_out0 = v_CIN_2365_out0[13:13];
assign v__8724_out0 = v_CIN_2380_out0[13:13];
assign v__8779_out0 = v_CIN_2365_out0[14:14];
assign v__8794_out0 = v_CIN_2380_out0[14:14];
assign v__10729_out0 = v_CIN_2365_out0[5:5];
assign v__10744_out0 = v_CIN_2380_out0[5:5];
assign v__13458_out0 = v_CIN_2365_out0[4:4];
assign v__13473_out0 = v_CIN_2380_out0[4:4];
assign v_RM_3504_out0 = v__7654_out0;
assign v_RM_3505_out0 = v__8779_out0;
assign v_RM_3507_out0 = v__10729_out0;
assign v_RM_3508_out0 = v__13458_out0;
assign v_RM_3509_out0 = v__8709_out0;
assign v_RM_3510_out0 = v__3061_out0;
assign v_RM_3511_out0 = v__3871_out0;
assign v_RM_3512_out0 = v__3833_out0;
assign v_RM_3513_out0 = v__2165_out0;
assign v_RM_3514_out0 = v__1783_out0;
assign v_RM_3515_out0 = v__3149_out0;
assign v_RM_3516_out0 = v__6810_out0;
assign v_RM_3517_out0 = v__478_out0;
assign v_RM_3518_out0 = v__3095_out0;
assign v_RM_3728_out0 = v__7669_out0;
assign v_RM_3729_out0 = v__8794_out0;
assign v_RM_3731_out0 = v__10744_out0;
assign v_RM_3732_out0 = v__13473_out0;
assign v_RM_3733_out0 = v__8724_out0;
assign v_RM_3734_out0 = v__3076_out0;
assign v_RM_3735_out0 = v__3886_out0;
assign v_RM_3736_out0 = v__3848_out0;
assign v_RM_3737_out0 = v__2180_out0;
assign v_RM_3738_out0 = v__1798_out0;
assign v_RM_3739_out0 = v__3164_out0;
assign v_RM_3740_out0 = v__6825_out0;
assign v_RM_3741_out0 = v__493_out0;
assign v_RM_3742_out0 = v__3110_out0;
assign v_CIN_9959_out0 = v__2204_out0;
assign v_CIN_10183_out0 = v__2218_out0;
assign v_RM_11623_out0 = v__2512_out0;
assign v_RM_12087_out0 = v__2527_out0;
assign v_RD_6176_out0 = v_CIN_9959_out0;
assign v_RD_6640_out0 = v_CIN_10183_out0;
assign v_G1_8038_out0 = ((v_RD_6183_out0 && !v_RM_11623_out0) || (!v_RD_6183_out0) && v_RM_11623_out0);
assign v_G1_8502_out0 = ((v_RD_6647_out0 && !v_RM_12087_out0) || (!v_RD_6647_out0) && v_RM_12087_out0);
assign v_RM_11611_out0 = v_RM_3504_out0;
assign v_RM_11613_out0 = v_RM_3505_out0;
assign v_RM_11617_out0 = v_RM_3507_out0;
assign v_RM_11619_out0 = v_RM_3508_out0;
assign v_RM_11621_out0 = v_RM_3509_out0;
assign v_RM_11624_out0 = v_RM_3510_out0;
assign v_RM_11626_out0 = v_RM_3511_out0;
assign v_RM_11628_out0 = v_RM_3512_out0;
assign v_RM_11630_out0 = v_RM_3513_out0;
assign v_RM_11632_out0 = v_RM_3514_out0;
assign v_RM_11634_out0 = v_RM_3515_out0;
assign v_RM_11636_out0 = v_RM_3516_out0;
assign v_RM_11638_out0 = v_RM_3517_out0;
assign v_RM_11640_out0 = v_RM_3518_out0;
assign v_RM_12075_out0 = v_RM_3728_out0;
assign v_RM_12077_out0 = v_RM_3729_out0;
assign v_RM_12081_out0 = v_RM_3731_out0;
assign v_RM_12083_out0 = v_RM_3732_out0;
assign v_RM_12085_out0 = v_RM_3733_out0;
assign v_RM_12088_out0 = v_RM_3734_out0;
assign v_RM_12090_out0 = v_RM_3735_out0;
assign v_RM_12092_out0 = v_RM_3736_out0;
assign v_RM_12094_out0 = v_RM_3737_out0;
assign v_RM_12096_out0 = v_RM_3738_out0;
assign v_RM_12098_out0 = v_RM_3739_out0;
assign v_RM_12100_out0 = v_RM_3740_out0;
assign v_RM_12102_out0 = v_RM_3741_out0;
assign v_RM_12104_out0 = v_RM_3742_out0;
assign v_G2_12574_out0 = v_RD_6183_out0 && v_RM_11623_out0;
assign v_G2_13038_out0 = v_RD_6647_out0 && v_RM_12087_out0;
assign v_CARRY_5183_out0 = v_G2_12574_out0;
assign v_CARRY_5647_out0 = v_G2_13038_out0;
assign v_G1_8026_out0 = ((v_RD_6171_out0 && !v_RM_11611_out0) || (!v_RD_6171_out0) && v_RM_11611_out0);
assign v_G1_8028_out0 = ((v_RD_6173_out0 && !v_RM_11613_out0) || (!v_RD_6173_out0) && v_RM_11613_out0);
assign v_G1_8032_out0 = ((v_RD_6177_out0 && !v_RM_11617_out0) || (!v_RD_6177_out0) && v_RM_11617_out0);
assign v_G1_8034_out0 = ((v_RD_6179_out0 && !v_RM_11619_out0) || (!v_RD_6179_out0) && v_RM_11619_out0);
assign v_G1_8036_out0 = ((v_RD_6181_out0 && !v_RM_11621_out0) || (!v_RD_6181_out0) && v_RM_11621_out0);
assign v_G1_8039_out0 = ((v_RD_6184_out0 && !v_RM_11624_out0) || (!v_RD_6184_out0) && v_RM_11624_out0);
assign v_G1_8041_out0 = ((v_RD_6186_out0 && !v_RM_11626_out0) || (!v_RD_6186_out0) && v_RM_11626_out0);
assign v_G1_8043_out0 = ((v_RD_6188_out0 && !v_RM_11628_out0) || (!v_RD_6188_out0) && v_RM_11628_out0);
assign v_G1_8045_out0 = ((v_RD_6190_out0 && !v_RM_11630_out0) || (!v_RD_6190_out0) && v_RM_11630_out0);
assign v_G1_8047_out0 = ((v_RD_6192_out0 && !v_RM_11632_out0) || (!v_RD_6192_out0) && v_RM_11632_out0);
assign v_G1_8049_out0 = ((v_RD_6194_out0 && !v_RM_11634_out0) || (!v_RD_6194_out0) && v_RM_11634_out0);
assign v_G1_8051_out0 = ((v_RD_6196_out0 && !v_RM_11636_out0) || (!v_RD_6196_out0) && v_RM_11636_out0);
assign v_G1_8053_out0 = ((v_RD_6198_out0 && !v_RM_11638_out0) || (!v_RD_6198_out0) && v_RM_11638_out0);
assign v_G1_8055_out0 = ((v_RD_6200_out0 && !v_RM_11640_out0) || (!v_RD_6200_out0) && v_RM_11640_out0);
assign v_G1_8490_out0 = ((v_RD_6635_out0 && !v_RM_12075_out0) || (!v_RD_6635_out0) && v_RM_12075_out0);
assign v_G1_8492_out0 = ((v_RD_6637_out0 && !v_RM_12077_out0) || (!v_RD_6637_out0) && v_RM_12077_out0);
assign v_G1_8496_out0 = ((v_RD_6641_out0 && !v_RM_12081_out0) || (!v_RD_6641_out0) && v_RM_12081_out0);
assign v_G1_8498_out0 = ((v_RD_6643_out0 && !v_RM_12083_out0) || (!v_RD_6643_out0) && v_RM_12083_out0);
assign v_G1_8500_out0 = ((v_RD_6645_out0 && !v_RM_12085_out0) || (!v_RD_6645_out0) && v_RM_12085_out0);
assign v_G1_8503_out0 = ((v_RD_6648_out0 && !v_RM_12088_out0) || (!v_RD_6648_out0) && v_RM_12088_out0);
assign v_G1_8505_out0 = ((v_RD_6650_out0 && !v_RM_12090_out0) || (!v_RD_6650_out0) && v_RM_12090_out0);
assign v_G1_8507_out0 = ((v_RD_6652_out0 && !v_RM_12092_out0) || (!v_RD_6652_out0) && v_RM_12092_out0);
assign v_G1_8509_out0 = ((v_RD_6654_out0 && !v_RM_12094_out0) || (!v_RD_6654_out0) && v_RM_12094_out0);
assign v_G1_8511_out0 = ((v_RD_6656_out0 && !v_RM_12096_out0) || (!v_RD_6656_out0) && v_RM_12096_out0);
assign v_G1_8513_out0 = ((v_RD_6658_out0 && !v_RM_12098_out0) || (!v_RD_6658_out0) && v_RM_12098_out0);
assign v_G1_8515_out0 = ((v_RD_6660_out0 && !v_RM_12100_out0) || (!v_RD_6660_out0) && v_RM_12100_out0);
assign v_G1_8517_out0 = ((v_RD_6662_out0 && !v_RM_12102_out0) || (!v_RD_6662_out0) && v_RM_12102_out0);
assign v_G1_8519_out0 = ((v_RD_6664_out0 && !v_RM_12104_out0) || (!v_RD_6664_out0) && v_RM_12104_out0);
assign v_S_9184_out0 = v_G1_8038_out0;
assign v_S_9648_out0 = v_G1_8502_out0;
assign v_G2_12562_out0 = v_RD_6171_out0 && v_RM_11611_out0;
assign v_G2_12564_out0 = v_RD_6173_out0 && v_RM_11613_out0;
assign v_G2_12568_out0 = v_RD_6177_out0 && v_RM_11617_out0;
assign v_G2_12570_out0 = v_RD_6179_out0 && v_RM_11619_out0;
assign v_G2_12572_out0 = v_RD_6181_out0 && v_RM_11621_out0;
assign v_G2_12575_out0 = v_RD_6184_out0 && v_RM_11624_out0;
assign v_G2_12577_out0 = v_RD_6186_out0 && v_RM_11626_out0;
assign v_G2_12579_out0 = v_RD_6188_out0 && v_RM_11628_out0;
assign v_G2_12581_out0 = v_RD_6190_out0 && v_RM_11630_out0;
assign v_G2_12583_out0 = v_RD_6192_out0 && v_RM_11632_out0;
assign v_G2_12585_out0 = v_RD_6194_out0 && v_RM_11634_out0;
assign v_G2_12587_out0 = v_RD_6196_out0 && v_RM_11636_out0;
assign v_G2_12589_out0 = v_RD_6198_out0 && v_RM_11638_out0;
assign v_G2_12591_out0 = v_RD_6200_out0 && v_RM_11640_out0;
assign v_G2_13026_out0 = v_RD_6635_out0 && v_RM_12075_out0;
assign v_G2_13028_out0 = v_RD_6637_out0 && v_RM_12077_out0;
assign v_G2_13032_out0 = v_RD_6641_out0 && v_RM_12081_out0;
assign v_G2_13034_out0 = v_RD_6643_out0 && v_RM_12083_out0;
assign v_G2_13036_out0 = v_RD_6645_out0 && v_RM_12085_out0;
assign v_G2_13039_out0 = v_RD_6648_out0 && v_RM_12088_out0;
assign v_G2_13041_out0 = v_RD_6650_out0 && v_RM_12090_out0;
assign v_G2_13043_out0 = v_RD_6652_out0 && v_RM_12092_out0;
assign v_G2_13045_out0 = v_RD_6654_out0 && v_RM_12094_out0;
assign v_G2_13047_out0 = v_RD_6656_out0 && v_RM_12096_out0;
assign v_G2_13049_out0 = v_RD_6658_out0 && v_RM_12098_out0;
assign v_G2_13051_out0 = v_RD_6660_out0 && v_RM_12100_out0;
assign v_G2_13053_out0 = v_RD_6662_out0 && v_RM_12102_out0;
assign v_G2_13055_out0 = v_RD_6664_out0 && v_RM_12104_out0;
assign v_S_4675_out0 = v_S_9184_out0;
assign v_S_4690_out0 = v_S_9648_out0;
assign v_CARRY_5171_out0 = v_G2_12562_out0;
assign v_CARRY_5173_out0 = v_G2_12564_out0;
assign v_CARRY_5177_out0 = v_G2_12568_out0;
assign v_CARRY_5179_out0 = v_G2_12570_out0;
assign v_CARRY_5181_out0 = v_G2_12572_out0;
assign v_CARRY_5184_out0 = v_G2_12575_out0;
assign v_CARRY_5186_out0 = v_G2_12577_out0;
assign v_CARRY_5188_out0 = v_G2_12579_out0;
assign v_CARRY_5190_out0 = v_G2_12581_out0;
assign v_CARRY_5192_out0 = v_G2_12583_out0;
assign v_CARRY_5194_out0 = v_G2_12585_out0;
assign v_CARRY_5196_out0 = v_G2_12587_out0;
assign v_CARRY_5198_out0 = v_G2_12589_out0;
assign v_CARRY_5200_out0 = v_G2_12591_out0;
assign v_CARRY_5635_out0 = v_G2_13026_out0;
assign v_CARRY_5637_out0 = v_G2_13028_out0;
assign v_CARRY_5641_out0 = v_G2_13032_out0;
assign v_CARRY_5643_out0 = v_G2_13034_out0;
assign v_CARRY_5645_out0 = v_G2_13036_out0;
assign v_CARRY_5648_out0 = v_G2_13039_out0;
assign v_CARRY_5650_out0 = v_G2_13041_out0;
assign v_CARRY_5652_out0 = v_G2_13043_out0;
assign v_CARRY_5654_out0 = v_G2_13045_out0;
assign v_CARRY_5656_out0 = v_G2_13047_out0;
assign v_CARRY_5658_out0 = v_G2_13049_out0;
assign v_CARRY_5660_out0 = v_G2_13051_out0;
assign v_CARRY_5662_out0 = v_G2_13053_out0;
assign v_CARRY_5664_out0 = v_G2_13055_out0;
assign v_S_9172_out0 = v_G1_8026_out0;
assign v_S_9174_out0 = v_G1_8028_out0;
assign v_S_9178_out0 = v_G1_8032_out0;
assign v_S_9180_out0 = v_G1_8034_out0;
assign v_S_9182_out0 = v_G1_8036_out0;
assign v_S_9185_out0 = v_G1_8039_out0;
assign v_S_9187_out0 = v_G1_8041_out0;
assign v_S_9189_out0 = v_G1_8043_out0;
assign v_S_9191_out0 = v_G1_8045_out0;
assign v_S_9193_out0 = v_G1_8047_out0;
assign v_S_9195_out0 = v_G1_8049_out0;
assign v_S_9197_out0 = v_G1_8051_out0;
assign v_S_9199_out0 = v_G1_8053_out0;
assign v_S_9201_out0 = v_G1_8055_out0;
assign v_S_9636_out0 = v_G1_8490_out0;
assign v_S_9638_out0 = v_G1_8492_out0;
assign v_S_9642_out0 = v_G1_8496_out0;
assign v_S_9644_out0 = v_G1_8498_out0;
assign v_S_9646_out0 = v_G1_8500_out0;
assign v_S_9649_out0 = v_G1_8503_out0;
assign v_S_9651_out0 = v_G1_8505_out0;
assign v_S_9653_out0 = v_G1_8507_out0;
assign v_S_9655_out0 = v_G1_8509_out0;
assign v_S_9657_out0 = v_G1_8511_out0;
assign v_S_9659_out0 = v_G1_8513_out0;
assign v_S_9661_out0 = v_G1_8515_out0;
assign v_S_9663_out0 = v_G1_8517_out0;
assign v_S_9665_out0 = v_G1_8519_out0;
assign v_CIN_9965_out0 = v_CARRY_5183_out0;
assign v_CIN_10189_out0 = v_CARRY_5647_out0;
assign v__56_out0 = { v__2392_out0,v_S_4675_out0 };
assign v__57_out0 = { v__2393_out0,v_S_4690_out0 };
assign v_RD_6189_out0 = v_CIN_9965_out0;
assign v_RD_6653_out0 = v_CIN_10189_out0;
assign v_RM_11612_out0 = v_S_9172_out0;
assign v_RM_11614_out0 = v_S_9174_out0;
assign v_RM_11618_out0 = v_S_9178_out0;
assign v_RM_11620_out0 = v_S_9180_out0;
assign v_RM_11622_out0 = v_S_9182_out0;
assign v_RM_11625_out0 = v_S_9185_out0;
assign v_RM_11627_out0 = v_S_9187_out0;
assign v_RM_11629_out0 = v_S_9189_out0;
assign v_RM_11631_out0 = v_S_9191_out0;
assign v_RM_11633_out0 = v_S_9193_out0;
assign v_RM_11635_out0 = v_S_9195_out0;
assign v_RM_11637_out0 = v_S_9197_out0;
assign v_RM_11639_out0 = v_S_9199_out0;
assign v_RM_11641_out0 = v_S_9201_out0;
assign v_RM_12076_out0 = v_S_9636_out0;
assign v_RM_12078_out0 = v_S_9638_out0;
assign v_RM_12082_out0 = v_S_9642_out0;
assign v_RM_12084_out0 = v_S_9644_out0;
assign v_RM_12086_out0 = v_S_9646_out0;
assign v_RM_12089_out0 = v_S_9649_out0;
assign v_RM_12091_out0 = v_S_9651_out0;
assign v_RM_12093_out0 = v_S_9653_out0;
assign v_RM_12095_out0 = v_S_9655_out0;
assign v_RM_12097_out0 = v_S_9657_out0;
assign v_RM_12099_out0 = v_S_9659_out0;
assign v_RM_12101_out0 = v_S_9661_out0;
assign v_RM_12103_out0 = v_S_9663_out0;
assign v_RM_12105_out0 = v_S_9665_out0;
assign v_G1_8044_out0 = ((v_RD_6189_out0 && !v_RM_11629_out0) || (!v_RD_6189_out0) && v_RM_11629_out0);
assign v_G1_8508_out0 = ((v_RD_6653_out0 && !v_RM_12093_out0) || (!v_RD_6653_out0) && v_RM_12093_out0);
assign v_G2_12580_out0 = v_RD_6189_out0 && v_RM_11629_out0;
assign v_G2_13044_out0 = v_RD_6653_out0 && v_RM_12093_out0;
assign v_CARRY_5189_out0 = v_G2_12580_out0;
assign v_CARRY_5653_out0 = v_G2_13044_out0;
assign v_S_9190_out0 = v_G1_8044_out0;
assign v_S_9654_out0 = v_G1_8508_out0;
assign v_S_1376_out0 = v_S_9190_out0;
assign v_S_1600_out0 = v_S_9654_out0;
assign v_G1_4152_out0 = v_CARRY_5189_out0 || v_CARRY_5188_out0;
assign v_G1_4376_out0 = v_CARRY_5653_out0 || v_CARRY_5652_out0;
assign v_COUT_844_out0 = v_G1_4152_out0;
assign v_COUT_1068_out0 = v_G1_4376_out0;
assign v_CIN_9971_out0 = v_COUT_844_out0;
assign v_CIN_10195_out0 = v_COUT_1068_out0;
assign v_RD_6201_out0 = v_CIN_9971_out0;
assign v_RD_6665_out0 = v_CIN_10195_out0;
assign v_G1_8056_out0 = ((v_RD_6201_out0 && !v_RM_11641_out0) || (!v_RD_6201_out0) && v_RM_11641_out0);
assign v_G1_8520_out0 = ((v_RD_6665_out0 && !v_RM_12105_out0) || (!v_RD_6665_out0) && v_RM_12105_out0);
assign v_G2_12592_out0 = v_RD_6201_out0 && v_RM_11641_out0;
assign v_G2_13056_out0 = v_RD_6665_out0 && v_RM_12105_out0;
assign v_CARRY_5201_out0 = v_G2_12592_out0;
assign v_CARRY_5665_out0 = v_G2_13056_out0;
assign v_S_9202_out0 = v_G1_8056_out0;
assign v_S_9666_out0 = v_G1_8520_out0;
assign v_S_1382_out0 = v_S_9202_out0;
assign v_S_1606_out0 = v_S_9666_out0;
assign v_G1_4158_out0 = v_CARRY_5201_out0 || v_CARRY_5200_out0;
assign v_G1_4382_out0 = v_CARRY_5665_out0 || v_CARRY_5664_out0;
assign v_COUT_850_out0 = v_G1_4158_out0;
assign v_COUT_1074_out0 = v_G1_4382_out0;
assign v__4792_out0 = { v_S_1376_out0,v_S_1382_out0 };
assign v__4807_out0 = { v_S_1600_out0,v_S_1606_out0 };
assign v_CIN_9966_out0 = v_COUT_850_out0;
assign v_CIN_10190_out0 = v_COUT_1074_out0;
assign v_RD_6191_out0 = v_CIN_9966_out0;
assign v_RD_6655_out0 = v_CIN_10190_out0;
assign v_G1_8046_out0 = ((v_RD_6191_out0 && !v_RM_11631_out0) || (!v_RD_6191_out0) && v_RM_11631_out0);
assign v_G1_8510_out0 = ((v_RD_6655_out0 && !v_RM_12095_out0) || (!v_RD_6655_out0) && v_RM_12095_out0);
assign v_G2_12582_out0 = v_RD_6191_out0 && v_RM_11631_out0;
assign v_G2_13046_out0 = v_RD_6655_out0 && v_RM_12095_out0;
assign v_CARRY_5191_out0 = v_G2_12582_out0;
assign v_CARRY_5655_out0 = v_G2_13046_out0;
assign v_S_9192_out0 = v_G1_8046_out0;
assign v_S_9656_out0 = v_G1_8510_out0;
assign v_S_1377_out0 = v_S_9192_out0;
assign v_S_1601_out0 = v_S_9656_out0;
assign v_G1_4153_out0 = v_CARRY_5191_out0 || v_CARRY_5190_out0;
assign v_G1_4377_out0 = v_CARRY_5655_out0 || v_CARRY_5654_out0;
assign v_COUT_845_out0 = v_G1_4153_out0;
assign v_COUT_1069_out0 = v_G1_4377_out0;
assign v__2562_out0 = { v__4792_out0,v_S_1377_out0 };
assign v__2577_out0 = { v__4807_out0,v_S_1601_out0 };
assign v_CIN_9961_out0 = v_COUT_845_out0;
assign v_CIN_10185_out0 = v_COUT_1069_out0;
assign v_RD_6180_out0 = v_CIN_9961_out0;
assign v_RD_6644_out0 = v_CIN_10185_out0;
assign v_G1_8035_out0 = ((v_RD_6180_out0 && !v_RM_11620_out0) || (!v_RD_6180_out0) && v_RM_11620_out0);
assign v_G1_8499_out0 = ((v_RD_6644_out0 && !v_RM_12084_out0) || (!v_RD_6644_out0) && v_RM_12084_out0);
assign v_G2_12571_out0 = v_RD_6180_out0 && v_RM_11620_out0;
assign v_G2_13035_out0 = v_RD_6644_out0 && v_RM_12084_out0;
assign v_CARRY_5180_out0 = v_G2_12571_out0;
assign v_CARRY_5644_out0 = v_G2_13035_out0;
assign v_S_9181_out0 = v_G1_8035_out0;
assign v_S_9645_out0 = v_G1_8499_out0;
assign v_S_1372_out0 = v_S_9181_out0;
assign v_S_1596_out0 = v_S_9645_out0;
assign v_G1_4148_out0 = v_CARRY_5180_out0 || v_CARRY_5179_out0;
assign v_G1_4372_out0 = v_CARRY_5644_out0 || v_CARRY_5643_out0;
assign v_COUT_840_out0 = v_G1_4148_out0;
assign v_COUT_1064_out0 = v_G1_4372_out0;
assign v__7042_out0 = { v__2562_out0,v_S_1372_out0 };
assign v__7057_out0 = { v__2577_out0,v_S_1596_out0 };
assign v_CIN_9960_out0 = v_COUT_840_out0;
assign v_CIN_10184_out0 = v_COUT_1064_out0;
assign v_RD_6178_out0 = v_CIN_9960_out0;
assign v_RD_6642_out0 = v_CIN_10184_out0;
assign v_G1_8033_out0 = ((v_RD_6178_out0 && !v_RM_11618_out0) || (!v_RD_6178_out0) && v_RM_11618_out0);
assign v_G1_8497_out0 = ((v_RD_6642_out0 && !v_RM_12082_out0) || (!v_RD_6642_out0) && v_RM_12082_out0);
assign v_G2_12569_out0 = v_RD_6178_out0 && v_RM_11618_out0;
assign v_G2_13033_out0 = v_RD_6642_out0 && v_RM_12082_out0;
assign v_CARRY_5178_out0 = v_G2_12569_out0;
assign v_CARRY_5642_out0 = v_G2_13033_out0;
assign v_S_9179_out0 = v_G1_8033_out0;
assign v_S_9643_out0 = v_G1_8497_out0;
assign v_S_1371_out0 = v_S_9179_out0;
assign v_S_1595_out0 = v_S_9643_out0;
assign v_G1_4147_out0 = v_CARRY_5178_out0 || v_CARRY_5177_out0;
assign v_G1_4371_out0 = v_CARRY_5642_out0 || v_CARRY_5641_out0;
assign v_COUT_839_out0 = v_G1_4147_out0;
assign v_COUT_1063_out0 = v_G1_4371_out0;
assign v__13528_out0 = { v__7042_out0,v_S_1371_out0 };
assign v__13543_out0 = { v__7057_out0,v_S_1595_out0 };
assign v_CIN_9967_out0 = v_COUT_839_out0;
assign v_CIN_10191_out0 = v_COUT_1063_out0;
assign v_RD_6193_out0 = v_CIN_9967_out0;
assign v_RD_6657_out0 = v_CIN_10191_out0;
assign v_G1_8048_out0 = ((v_RD_6193_out0 && !v_RM_11633_out0) || (!v_RD_6193_out0) && v_RM_11633_out0);
assign v_G1_8512_out0 = ((v_RD_6657_out0 && !v_RM_12097_out0) || (!v_RD_6657_out0) && v_RM_12097_out0);
assign v_G2_12584_out0 = v_RD_6193_out0 && v_RM_11633_out0;
assign v_G2_13048_out0 = v_RD_6657_out0 && v_RM_12097_out0;
assign v_CARRY_5193_out0 = v_G2_12584_out0;
assign v_CARRY_5657_out0 = v_G2_13048_out0;
assign v_S_9194_out0 = v_G1_8048_out0;
assign v_S_9658_out0 = v_G1_8512_out0;
assign v_S_1378_out0 = v_S_9194_out0;
assign v_S_1602_out0 = v_S_9658_out0;
assign v_G1_4154_out0 = v_CARRY_5193_out0 || v_CARRY_5192_out0;
assign v_G1_4378_out0 = v_CARRY_5657_out0 || v_CARRY_5656_out0;
assign v_COUT_846_out0 = v_G1_4154_out0;
assign v_COUT_1070_out0 = v_G1_4378_out0;
assign v__3321_out0 = { v__13528_out0,v_S_1378_out0 };
assign v__3336_out0 = { v__13543_out0,v_S_1602_out0 };
assign v_CIN_9968_out0 = v_COUT_846_out0;
assign v_CIN_10192_out0 = v_COUT_1070_out0;
assign v_RD_6195_out0 = v_CIN_9968_out0;
assign v_RD_6659_out0 = v_CIN_10192_out0;
assign v_G1_8050_out0 = ((v_RD_6195_out0 && !v_RM_11635_out0) || (!v_RD_6195_out0) && v_RM_11635_out0);
assign v_G1_8514_out0 = ((v_RD_6659_out0 && !v_RM_12099_out0) || (!v_RD_6659_out0) && v_RM_12099_out0);
assign v_G2_12586_out0 = v_RD_6195_out0 && v_RM_11635_out0;
assign v_G2_13050_out0 = v_RD_6659_out0 && v_RM_12099_out0;
assign v_CARRY_5195_out0 = v_G2_12586_out0;
assign v_CARRY_5659_out0 = v_G2_13050_out0;
assign v_S_9196_out0 = v_G1_8050_out0;
assign v_S_9660_out0 = v_G1_8514_out0;
assign v_S_1379_out0 = v_S_9196_out0;
assign v_S_1603_out0 = v_S_9660_out0;
assign v_G1_4155_out0 = v_CARRY_5195_out0 || v_CARRY_5194_out0;
assign v_G1_4379_out0 = v_CARRY_5659_out0 || v_CARRY_5658_out0;
assign v_COUT_847_out0 = v_G1_4155_out0;
assign v_COUT_1071_out0 = v_G1_4379_out0;
assign v__7157_out0 = { v__3321_out0,v_S_1379_out0 };
assign v__7172_out0 = { v__3336_out0,v_S_1603_out0 };
assign v_CIN_9970_out0 = v_COUT_847_out0;
assign v_CIN_10194_out0 = v_COUT_1071_out0;
assign v_RD_6199_out0 = v_CIN_9970_out0;
assign v_RD_6663_out0 = v_CIN_10194_out0;
assign v_G1_8054_out0 = ((v_RD_6199_out0 && !v_RM_11639_out0) || (!v_RD_6199_out0) && v_RM_11639_out0);
assign v_G1_8518_out0 = ((v_RD_6663_out0 && !v_RM_12103_out0) || (!v_RD_6663_out0) && v_RM_12103_out0);
assign v_G2_12590_out0 = v_RD_6199_out0 && v_RM_11639_out0;
assign v_G2_13054_out0 = v_RD_6663_out0 && v_RM_12103_out0;
assign v_CARRY_5199_out0 = v_G2_12590_out0;
assign v_CARRY_5663_out0 = v_G2_13054_out0;
assign v_S_9200_out0 = v_G1_8054_out0;
assign v_S_9664_out0 = v_G1_8518_out0;
assign v_S_1381_out0 = v_S_9200_out0;
assign v_S_1605_out0 = v_S_9664_out0;
assign v_G1_4157_out0 = v_CARRY_5199_out0 || v_CARRY_5198_out0;
assign v_G1_4381_out0 = v_CARRY_5663_out0 || v_CARRY_5662_out0;
assign v_COUT_849_out0 = v_G1_4157_out0;
assign v_COUT_1073_out0 = v_G1_4381_out0;
assign v__4759_out0 = { v__7157_out0,v_S_1381_out0 };
assign v__4774_out0 = { v__7172_out0,v_S_1605_out0 };
assign v_CIN_9963_out0 = v_COUT_849_out0;
assign v_CIN_10187_out0 = v_COUT_1073_out0;
assign v_RD_6185_out0 = v_CIN_9963_out0;
assign v_RD_6649_out0 = v_CIN_10187_out0;
assign v_G1_8040_out0 = ((v_RD_6185_out0 && !v_RM_11625_out0) || (!v_RD_6185_out0) && v_RM_11625_out0);
assign v_G1_8504_out0 = ((v_RD_6649_out0 && !v_RM_12089_out0) || (!v_RD_6649_out0) && v_RM_12089_out0);
assign v_G2_12576_out0 = v_RD_6185_out0 && v_RM_11625_out0;
assign v_G2_13040_out0 = v_RD_6649_out0 && v_RM_12089_out0;
assign v_CARRY_5185_out0 = v_G2_12576_out0;
assign v_CARRY_5649_out0 = v_G2_13040_out0;
assign v_S_9186_out0 = v_G1_8040_out0;
assign v_S_9650_out0 = v_G1_8504_out0;
assign v_S_1374_out0 = v_S_9186_out0;
assign v_S_1598_out0 = v_S_9650_out0;
assign v_G1_4150_out0 = v_CARRY_5185_out0 || v_CARRY_5184_out0;
assign v_G1_4374_out0 = v_CARRY_5649_out0 || v_CARRY_5648_out0;
assign v_COUT_842_out0 = v_G1_4150_out0;
assign v_COUT_1066_out0 = v_G1_4374_out0;
assign v__6936_out0 = { v__4759_out0,v_S_1374_out0 };
assign v__6951_out0 = { v__4774_out0,v_S_1598_out0 };
assign v_CIN_9964_out0 = v_COUT_842_out0;
assign v_CIN_10188_out0 = v_COUT_1066_out0;
assign v_RD_6187_out0 = v_CIN_9964_out0;
assign v_RD_6651_out0 = v_CIN_10188_out0;
assign v_G1_8042_out0 = ((v_RD_6187_out0 && !v_RM_11627_out0) || (!v_RD_6187_out0) && v_RM_11627_out0);
assign v_G1_8506_out0 = ((v_RD_6651_out0 && !v_RM_12091_out0) || (!v_RD_6651_out0) && v_RM_12091_out0);
assign v_G2_12578_out0 = v_RD_6187_out0 && v_RM_11627_out0;
assign v_G2_13042_out0 = v_RD_6651_out0 && v_RM_12091_out0;
assign v_CARRY_5187_out0 = v_G2_12578_out0;
assign v_CARRY_5651_out0 = v_G2_13042_out0;
assign v_S_9188_out0 = v_G1_8042_out0;
assign v_S_9652_out0 = v_G1_8506_out0;
assign v_S_1375_out0 = v_S_9188_out0;
assign v_S_1599_out0 = v_S_9652_out0;
assign v_G1_4151_out0 = v_CARRY_5187_out0 || v_CARRY_5186_out0;
assign v_G1_4375_out0 = v_CARRY_5651_out0 || v_CARRY_5650_out0;
assign v_COUT_843_out0 = v_G1_4151_out0;
assign v_COUT_1067_out0 = v_G1_4375_out0;
assign v__5812_out0 = { v__6936_out0,v_S_1375_out0 };
assign v__5827_out0 = { v__6951_out0,v_S_1599_out0 };
assign v_CIN_9969_out0 = v_COUT_843_out0;
assign v_CIN_10193_out0 = v_COUT_1067_out0;
assign v_RD_6197_out0 = v_CIN_9969_out0;
assign v_RD_6661_out0 = v_CIN_10193_out0;
assign v_G1_8052_out0 = ((v_RD_6197_out0 && !v_RM_11637_out0) || (!v_RD_6197_out0) && v_RM_11637_out0);
assign v_G1_8516_out0 = ((v_RD_6661_out0 && !v_RM_12101_out0) || (!v_RD_6661_out0) && v_RM_12101_out0);
assign v_G2_12588_out0 = v_RD_6197_out0 && v_RM_11637_out0;
assign v_G2_13052_out0 = v_RD_6661_out0 && v_RM_12101_out0;
assign v_CARRY_5197_out0 = v_G2_12588_out0;
assign v_CARRY_5661_out0 = v_G2_13052_out0;
assign v_S_9198_out0 = v_G1_8052_out0;
assign v_S_9662_out0 = v_G1_8516_out0;
assign v_S_1380_out0 = v_S_9198_out0;
assign v_S_1604_out0 = v_S_9662_out0;
assign v_G1_4156_out0 = v_CARRY_5197_out0 || v_CARRY_5196_out0;
assign v_G1_4380_out0 = v_CARRY_5661_out0 || v_CARRY_5660_out0;
assign v_COUT_848_out0 = v_G1_4156_out0;
assign v_COUT_1072_out0 = v_G1_4380_out0;
assign v__2036_out0 = { v__5812_out0,v_S_1380_out0 };
assign v__2051_out0 = { v__5827_out0,v_S_1604_out0 };
assign v_CIN_9957_out0 = v_COUT_848_out0;
assign v_CIN_10181_out0 = v_COUT_1072_out0;
assign v_RD_6172_out0 = v_CIN_9957_out0;
assign v_RD_6636_out0 = v_CIN_10181_out0;
assign v_G1_8027_out0 = ((v_RD_6172_out0 && !v_RM_11612_out0) || (!v_RD_6172_out0) && v_RM_11612_out0);
assign v_G1_8491_out0 = ((v_RD_6636_out0 && !v_RM_12076_out0) || (!v_RD_6636_out0) && v_RM_12076_out0);
assign v_G2_12563_out0 = v_RD_6172_out0 && v_RM_11612_out0;
assign v_G2_13027_out0 = v_RD_6636_out0 && v_RM_12076_out0;
assign v_CARRY_5172_out0 = v_G2_12563_out0;
assign v_CARRY_5636_out0 = v_G2_13027_out0;
assign v_S_9173_out0 = v_G1_8027_out0;
assign v_S_9637_out0 = v_G1_8491_out0;
assign v_S_1368_out0 = v_S_9173_out0;
assign v_S_1592_out0 = v_S_9637_out0;
assign v_G1_4144_out0 = v_CARRY_5172_out0 || v_CARRY_5171_out0;
assign v_G1_4368_out0 = v_CARRY_5636_out0 || v_CARRY_5635_out0;
assign v_COUT_836_out0 = v_G1_4144_out0;
assign v_COUT_1060_out0 = v_G1_4368_out0;
assign v__2803_out0 = { v__2036_out0,v_S_1368_out0 };
assign v__2818_out0 = { v__2051_out0,v_S_1592_out0 };
assign v_CIN_9962_out0 = v_COUT_836_out0;
assign v_CIN_10186_out0 = v_COUT_1060_out0;
assign v_RD_6182_out0 = v_CIN_9962_out0;
assign v_RD_6646_out0 = v_CIN_10186_out0;
assign v_G1_8037_out0 = ((v_RD_6182_out0 && !v_RM_11622_out0) || (!v_RD_6182_out0) && v_RM_11622_out0);
assign v_G1_8501_out0 = ((v_RD_6646_out0 && !v_RM_12086_out0) || (!v_RD_6646_out0) && v_RM_12086_out0);
assign v_G2_12573_out0 = v_RD_6182_out0 && v_RM_11622_out0;
assign v_G2_13037_out0 = v_RD_6646_out0 && v_RM_12086_out0;
assign v_CARRY_5182_out0 = v_G2_12573_out0;
assign v_CARRY_5646_out0 = v_G2_13037_out0;
assign v_S_9183_out0 = v_G1_8037_out0;
assign v_S_9647_out0 = v_G1_8501_out0;
assign v_S_1373_out0 = v_S_9183_out0;
assign v_S_1597_out0 = v_S_9647_out0;
assign v_G1_4149_out0 = v_CARRY_5182_out0 || v_CARRY_5181_out0;
assign v_G1_4373_out0 = v_CARRY_5646_out0 || v_CARRY_5645_out0;
assign v_COUT_841_out0 = v_G1_4149_out0;
assign v_COUT_1065_out0 = v_G1_4373_out0;
assign v__1835_out0 = { v__2803_out0,v_S_1373_out0 };
assign v__1850_out0 = { v__2818_out0,v_S_1597_out0 };
assign v_CIN_9958_out0 = v_COUT_841_out0;
assign v_CIN_10182_out0 = v_COUT_1065_out0;
assign v_RD_6174_out0 = v_CIN_9958_out0;
assign v_RD_6638_out0 = v_CIN_10182_out0;
assign v_G1_8029_out0 = ((v_RD_6174_out0 && !v_RM_11614_out0) || (!v_RD_6174_out0) && v_RM_11614_out0);
assign v_G1_8493_out0 = ((v_RD_6638_out0 && !v_RM_12078_out0) || (!v_RD_6638_out0) && v_RM_12078_out0);
assign v_G2_12565_out0 = v_RD_6174_out0 && v_RM_11614_out0;
assign v_G2_13029_out0 = v_RD_6638_out0 && v_RM_12078_out0;
assign v_CARRY_5174_out0 = v_G2_12565_out0;
assign v_CARRY_5638_out0 = v_G2_13029_out0;
assign v_S_9175_out0 = v_G1_8029_out0;
assign v_S_9639_out0 = v_G1_8493_out0;
assign v_S_1369_out0 = v_S_9175_out0;
assign v_S_1593_out0 = v_S_9639_out0;
assign v_G1_4145_out0 = v_CARRY_5174_out0 || v_CARRY_5173_out0;
assign v_G1_4369_out0 = v_CARRY_5638_out0 || v_CARRY_5637_out0;
assign v_COUT_837_out0 = v_G1_4145_out0;
assign v_COUT_1061_out0 = v_G1_4369_out0;
assign v__4559_out0 = { v__1835_out0,v_S_1369_out0 };
assign v__4574_out0 = { v__1850_out0,v_S_1593_out0 };
assign v_RM_3506_out0 = v_COUT_837_out0;
assign v_RM_3730_out0 = v_COUT_1061_out0;
assign v_RM_11615_out0 = v_RM_3506_out0;
assign v_RM_12079_out0 = v_RM_3730_out0;
assign v_G1_8030_out0 = ((v_RD_6175_out0 && !v_RM_11615_out0) || (!v_RD_6175_out0) && v_RM_11615_out0);
assign v_G1_8494_out0 = ((v_RD_6639_out0 && !v_RM_12079_out0) || (!v_RD_6639_out0) && v_RM_12079_out0);
assign v_G2_12566_out0 = v_RD_6175_out0 && v_RM_11615_out0;
assign v_G2_13030_out0 = v_RD_6639_out0 && v_RM_12079_out0;
assign v_CARRY_5175_out0 = v_G2_12566_out0;
assign v_CARRY_5639_out0 = v_G2_13030_out0;
assign v_S_9176_out0 = v_G1_8030_out0;
assign v_S_9640_out0 = v_G1_8494_out0;
assign v_RM_11616_out0 = v_S_9176_out0;
assign v_RM_12080_out0 = v_S_9640_out0;
assign v_G1_8031_out0 = ((v_RD_6176_out0 && !v_RM_11616_out0) || (!v_RD_6176_out0) && v_RM_11616_out0);
assign v_G1_8495_out0 = ((v_RD_6640_out0 && !v_RM_12080_out0) || (!v_RD_6640_out0) && v_RM_12080_out0);
assign v_G2_12567_out0 = v_RD_6176_out0 && v_RM_11616_out0;
assign v_G2_13031_out0 = v_RD_6640_out0 && v_RM_12080_out0;
assign v_CARRY_5176_out0 = v_G2_12567_out0;
assign v_CARRY_5640_out0 = v_G2_13031_out0;
assign v_S_9177_out0 = v_G1_8031_out0;
assign v_S_9641_out0 = v_G1_8495_out0;
assign v_S_1370_out0 = v_S_9177_out0;
assign v_S_1594_out0 = v_S_9641_out0;
assign v_G1_4146_out0 = v_CARRY_5176_out0 || v_CARRY_5175_out0;
assign v_G1_4370_out0 = v_CARRY_5640_out0 || v_CARRY_5639_out0;
assign v_COUT_838_out0 = v_G1_4146_out0;
assign v_COUT_1062_out0 = v_G1_4370_out0;
assign v__10661_out0 = { v__4559_out0,v_S_1370_out0 };
assign v__10676_out0 = { v__4574_out0,v_S_1594_out0 };
assign v__10956_out0 = { v__10661_out0,v_COUT_838_out0 };
assign v__10971_out0 = { v__10676_out0,v_COUT_1062_out0 };
assign v_COUT_10926_out0 = v__10956_out0;
assign v_COUT_10941_out0 = v__10971_out0;
assign v_CIN_2368_out0 = v_COUT_10926_out0;
assign v_CIN_2383_out0 = v_COUT_10941_out0;
assign v__481_out0 = v_CIN_2368_out0[8:8];
assign v__496_out0 = v_CIN_2383_out0[8:8];
assign v__1786_out0 = v_CIN_2368_out0[6:6];
assign v__1801_out0 = v_CIN_2383_out0[6:6];
assign v__2168_out0 = v_CIN_2368_out0[3:3];
assign v__2183_out0 = v_CIN_2383_out0[3:3];
assign v__2207_out0 = v_CIN_2368_out0[15:15];
assign v__2221_out0 = v_CIN_2383_out0[15:15];
assign v__2515_out0 = v_CIN_2368_out0[0:0];
assign v__2530_out0 = v_CIN_2383_out0[0:0];
assign v__3064_out0 = v_CIN_2368_out0[9:9];
assign v__3079_out0 = v_CIN_2383_out0[9:9];
assign v__3098_out0 = v_CIN_2368_out0[2:2];
assign v__3113_out0 = v_CIN_2383_out0[2:2];
assign v__3152_out0 = v_CIN_2368_out0[7:7];
assign v__3167_out0 = v_CIN_2383_out0[7:7];
assign v__3836_out0 = v_CIN_2368_out0[1:1];
assign v__3851_out0 = v_CIN_2383_out0[1:1];
assign v__3874_out0 = v_CIN_2368_out0[10:10];
assign v__3889_out0 = v_CIN_2383_out0[10:10];
assign v__6813_out0 = v_CIN_2368_out0[11:11];
assign v__6828_out0 = v_CIN_2383_out0[11:11];
assign v__7657_out0 = v_CIN_2368_out0[12:12];
assign v__7672_out0 = v_CIN_2383_out0[12:12];
assign v__8712_out0 = v_CIN_2368_out0[13:13];
assign v__8727_out0 = v_CIN_2383_out0[13:13];
assign v__8782_out0 = v_CIN_2368_out0[14:14];
assign v__8797_out0 = v_CIN_2383_out0[14:14];
assign v__10732_out0 = v_CIN_2368_out0[5:5];
assign v__10747_out0 = v_CIN_2383_out0[5:5];
assign v__13461_out0 = v_CIN_2368_out0[4:4];
assign v__13476_out0 = v_CIN_2383_out0[4:4];
assign v_RM_3549_out0 = v__7657_out0;
assign v_RM_3550_out0 = v__8782_out0;
assign v_RM_3552_out0 = v__10732_out0;
assign v_RM_3553_out0 = v__13461_out0;
assign v_RM_3554_out0 = v__8712_out0;
assign v_RM_3555_out0 = v__3064_out0;
assign v_RM_3556_out0 = v__3874_out0;
assign v_RM_3557_out0 = v__3836_out0;
assign v_RM_3558_out0 = v__2168_out0;
assign v_RM_3559_out0 = v__1786_out0;
assign v_RM_3560_out0 = v__3152_out0;
assign v_RM_3561_out0 = v__6813_out0;
assign v_RM_3562_out0 = v__481_out0;
assign v_RM_3563_out0 = v__3098_out0;
assign v_RM_3773_out0 = v__7672_out0;
assign v_RM_3774_out0 = v__8797_out0;
assign v_RM_3776_out0 = v__10747_out0;
assign v_RM_3777_out0 = v__13476_out0;
assign v_RM_3778_out0 = v__8727_out0;
assign v_RM_3779_out0 = v__3079_out0;
assign v_RM_3780_out0 = v__3889_out0;
assign v_RM_3781_out0 = v__3851_out0;
assign v_RM_3782_out0 = v__2183_out0;
assign v_RM_3783_out0 = v__1801_out0;
assign v_RM_3784_out0 = v__3167_out0;
assign v_RM_3785_out0 = v__6828_out0;
assign v_RM_3786_out0 = v__496_out0;
assign v_RM_3787_out0 = v__3113_out0;
assign v_CIN_10004_out0 = v__2207_out0;
assign v_CIN_10228_out0 = v__2221_out0;
assign v_RM_11716_out0 = v__2515_out0;
assign v_RM_12180_out0 = v__2530_out0;
assign v_RD_6269_out0 = v_CIN_10004_out0;
assign v_RD_6733_out0 = v_CIN_10228_out0;
assign v_G1_8131_out0 = ((v_RD_6276_out0 && !v_RM_11716_out0) || (!v_RD_6276_out0) && v_RM_11716_out0);
assign v_G1_8595_out0 = ((v_RD_6740_out0 && !v_RM_12180_out0) || (!v_RD_6740_out0) && v_RM_12180_out0);
assign v_RM_11704_out0 = v_RM_3549_out0;
assign v_RM_11706_out0 = v_RM_3550_out0;
assign v_RM_11710_out0 = v_RM_3552_out0;
assign v_RM_11712_out0 = v_RM_3553_out0;
assign v_RM_11714_out0 = v_RM_3554_out0;
assign v_RM_11717_out0 = v_RM_3555_out0;
assign v_RM_11719_out0 = v_RM_3556_out0;
assign v_RM_11721_out0 = v_RM_3557_out0;
assign v_RM_11723_out0 = v_RM_3558_out0;
assign v_RM_11725_out0 = v_RM_3559_out0;
assign v_RM_11727_out0 = v_RM_3560_out0;
assign v_RM_11729_out0 = v_RM_3561_out0;
assign v_RM_11731_out0 = v_RM_3562_out0;
assign v_RM_11733_out0 = v_RM_3563_out0;
assign v_RM_12168_out0 = v_RM_3773_out0;
assign v_RM_12170_out0 = v_RM_3774_out0;
assign v_RM_12174_out0 = v_RM_3776_out0;
assign v_RM_12176_out0 = v_RM_3777_out0;
assign v_RM_12178_out0 = v_RM_3778_out0;
assign v_RM_12181_out0 = v_RM_3779_out0;
assign v_RM_12183_out0 = v_RM_3780_out0;
assign v_RM_12185_out0 = v_RM_3781_out0;
assign v_RM_12187_out0 = v_RM_3782_out0;
assign v_RM_12189_out0 = v_RM_3783_out0;
assign v_RM_12191_out0 = v_RM_3784_out0;
assign v_RM_12193_out0 = v_RM_3785_out0;
assign v_RM_12195_out0 = v_RM_3786_out0;
assign v_RM_12197_out0 = v_RM_3787_out0;
assign v_G2_12667_out0 = v_RD_6276_out0 && v_RM_11716_out0;
assign v_G2_13131_out0 = v_RD_6740_out0 && v_RM_12180_out0;
assign v_CARRY_5276_out0 = v_G2_12667_out0;
assign v_CARRY_5740_out0 = v_G2_13131_out0;
assign v_G1_8119_out0 = ((v_RD_6264_out0 && !v_RM_11704_out0) || (!v_RD_6264_out0) && v_RM_11704_out0);
assign v_G1_8121_out0 = ((v_RD_6266_out0 && !v_RM_11706_out0) || (!v_RD_6266_out0) && v_RM_11706_out0);
assign v_G1_8125_out0 = ((v_RD_6270_out0 && !v_RM_11710_out0) || (!v_RD_6270_out0) && v_RM_11710_out0);
assign v_G1_8127_out0 = ((v_RD_6272_out0 && !v_RM_11712_out0) || (!v_RD_6272_out0) && v_RM_11712_out0);
assign v_G1_8129_out0 = ((v_RD_6274_out0 && !v_RM_11714_out0) || (!v_RD_6274_out0) && v_RM_11714_out0);
assign v_G1_8132_out0 = ((v_RD_6277_out0 && !v_RM_11717_out0) || (!v_RD_6277_out0) && v_RM_11717_out0);
assign v_G1_8134_out0 = ((v_RD_6279_out0 && !v_RM_11719_out0) || (!v_RD_6279_out0) && v_RM_11719_out0);
assign v_G1_8136_out0 = ((v_RD_6281_out0 && !v_RM_11721_out0) || (!v_RD_6281_out0) && v_RM_11721_out0);
assign v_G1_8138_out0 = ((v_RD_6283_out0 && !v_RM_11723_out0) || (!v_RD_6283_out0) && v_RM_11723_out0);
assign v_G1_8140_out0 = ((v_RD_6285_out0 && !v_RM_11725_out0) || (!v_RD_6285_out0) && v_RM_11725_out0);
assign v_G1_8142_out0 = ((v_RD_6287_out0 && !v_RM_11727_out0) || (!v_RD_6287_out0) && v_RM_11727_out0);
assign v_G1_8144_out0 = ((v_RD_6289_out0 && !v_RM_11729_out0) || (!v_RD_6289_out0) && v_RM_11729_out0);
assign v_G1_8146_out0 = ((v_RD_6291_out0 && !v_RM_11731_out0) || (!v_RD_6291_out0) && v_RM_11731_out0);
assign v_G1_8148_out0 = ((v_RD_6293_out0 && !v_RM_11733_out0) || (!v_RD_6293_out0) && v_RM_11733_out0);
assign v_G1_8583_out0 = ((v_RD_6728_out0 && !v_RM_12168_out0) || (!v_RD_6728_out0) && v_RM_12168_out0);
assign v_G1_8585_out0 = ((v_RD_6730_out0 && !v_RM_12170_out0) || (!v_RD_6730_out0) && v_RM_12170_out0);
assign v_G1_8589_out0 = ((v_RD_6734_out0 && !v_RM_12174_out0) || (!v_RD_6734_out0) && v_RM_12174_out0);
assign v_G1_8591_out0 = ((v_RD_6736_out0 && !v_RM_12176_out0) || (!v_RD_6736_out0) && v_RM_12176_out0);
assign v_G1_8593_out0 = ((v_RD_6738_out0 && !v_RM_12178_out0) || (!v_RD_6738_out0) && v_RM_12178_out0);
assign v_G1_8596_out0 = ((v_RD_6741_out0 && !v_RM_12181_out0) || (!v_RD_6741_out0) && v_RM_12181_out0);
assign v_G1_8598_out0 = ((v_RD_6743_out0 && !v_RM_12183_out0) || (!v_RD_6743_out0) && v_RM_12183_out0);
assign v_G1_8600_out0 = ((v_RD_6745_out0 && !v_RM_12185_out0) || (!v_RD_6745_out0) && v_RM_12185_out0);
assign v_G1_8602_out0 = ((v_RD_6747_out0 && !v_RM_12187_out0) || (!v_RD_6747_out0) && v_RM_12187_out0);
assign v_G1_8604_out0 = ((v_RD_6749_out0 && !v_RM_12189_out0) || (!v_RD_6749_out0) && v_RM_12189_out0);
assign v_G1_8606_out0 = ((v_RD_6751_out0 && !v_RM_12191_out0) || (!v_RD_6751_out0) && v_RM_12191_out0);
assign v_G1_8608_out0 = ((v_RD_6753_out0 && !v_RM_12193_out0) || (!v_RD_6753_out0) && v_RM_12193_out0);
assign v_G1_8610_out0 = ((v_RD_6755_out0 && !v_RM_12195_out0) || (!v_RD_6755_out0) && v_RM_12195_out0);
assign v_G1_8612_out0 = ((v_RD_6757_out0 && !v_RM_12197_out0) || (!v_RD_6757_out0) && v_RM_12197_out0);
assign v_S_9277_out0 = v_G1_8131_out0;
assign v_S_9741_out0 = v_G1_8595_out0;
assign v_G2_12655_out0 = v_RD_6264_out0 && v_RM_11704_out0;
assign v_G2_12657_out0 = v_RD_6266_out0 && v_RM_11706_out0;
assign v_G2_12661_out0 = v_RD_6270_out0 && v_RM_11710_out0;
assign v_G2_12663_out0 = v_RD_6272_out0 && v_RM_11712_out0;
assign v_G2_12665_out0 = v_RD_6274_out0 && v_RM_11714_out0;
assign v_G2_12668_out0 = v_RD_6277_out0 && v_RM_11717_out0;
assign v_G2_12670_out0 = v_RD_6279_out0 && v_RM_11719_out0;
assign v_G2_12672_out0 = v_RD_6281_out0 && v_RM_11721_out0;
assign v_G2_12674_out0 = v_RD_6283_out0 && v_RM_11723_out0;
assign v_G2_12676_out0 = v_RD_6285_out0 && v_RM_11725_out0;
assign v_G2_12678_out0 = v_RD_6287_out0 && v_RM_11727_out0;
assign v_G2_12680_out0 = v_RD_6289_out0 && v_RM_11729_out0;
assign v_G2_12682_out0 = v_RD_6291_out0 && v_RM_11731_out0;
assign v_G2_12684_out0 = v_RD_6293_out0 && v_RM_11733_out0;
assign v_G2_13119_out0 = v_RD_6728_out0 && v_RM_12168_out0;
assign v_G2_13121_out0 = v_RD_6730_out0 && v_RM_12170_out0;
assign v_G2_13125_out0 = v_RD_6734_out0 && v_RM_12174_out0;
assign v_G2_13127_out0 = v_RD_6736_out0 && v_RM_12176_out0;
assign v_G2_13129_out0 = v_RD_6738_out0 && v_RM_12178_out0;
assign v_G2_13132_out0 = v_RD_6741_out0 && v_RM_12181_out0;
assign v_G2_13134_out0 = v_RD_6743_out0 && v_RM_12183_out0;
assign v_G2_13136_out0 = v_RD_6745_out0 && v_RM_12185_out0;
assign v_G2_13138_out0 = v_RD_6747_out0 && v_RM_12187_out0;
assign v_G2_13140_out0 = v_RD_6749_out0 && v_RM_12189_out0;
assign v_G2_13142_out0 = v_RD_6751_out0 && v_RM_12191_out0;
assign v_G2_13144_out0 = v_RD_6753_out0 && v_RM_12193_out0;
assign v_G2_13146_out0 = v_RD_6755_out0 && v_RM_12195_out0;
assign v_G2_13148_out0 = v_RD_6757_out0 && v_RM_12197_out0;
assign v_S_4678_out0 = v_S_9277_out0;
assign v_S_4693_out0 = v_S_9741_out0;
assign v_CARRY_5264_out0 = v_G2_12655_out0;
assign v_CARRY_5266_out0 = v_G2_12657_out0;
assign v_CARRY_5270_out0 = v_G2_12661_out0;
assign v_CARRY_5272_out0 = v_G2_12663_out0;
assign v_CARRY_5274_out0 = v_G2_12665_out0;
assign v_CARRY_5277_out0 = v_G2_12668_out0;
assign v_CARRY_5279_out0 = v_G2_12670_out0;
assign v_CARRY_5281_out0 = v_G2_12672_out0;
assign v_CARRY_5283_out0 = v_G2_12674_out0;
assign v_CARRY_5285_out0 = v_G2_12676_out0;
assign v_CARRY_5287_out0 = v_G2_12678_out0;
assign v_CARRY_5289_out0 = v_G2_12680_out0;
assign v_CARRY_5291_out0 = v_G2_12682_out0;
assign v_CARRY_5293_out0 = v_G2_12684_out0;
assign v_CARRY_5728_out0 = v_G2_13119_out0;
assign v_CARRY_5730_out0 = v_G2_13121_out0;
assign v_CARRY_5734_out0 = v_G2_13125_out0;
assign v_CARRY_5736_out0 = v_G2_13127_out0;
assign v_CARRY_5738_out0 = v_G2_13129_out0;
assign v_CARRY_5741_out0 = v_G2_13132_out0;
assign v_CARRY_5743_out0 = v_G2_13134_out0;
assign v_CARRY_5745_out0 = v_G2_13136_out0;
assign v_CARRY_5747_out0 = v_G2_13138_out0;
assign v_CARRY_5749_out0 = v_G2_13140_out0;
assign v_CARRY_5751_out0 = v_G2_13142_out0;
assign v_CARRY_5753_out0 = v_G2_13144_out0;
assign v_CARRY_5755_out0 = v_G2_13146_out0;
assign v_CARRY_5757_out0 = v_G2_13148_out0;
assign v_S_9265_out0 = v_G1_8119_out0;
assign v_S_9267_out0 = v_G1_8121_out0;
assign v_S_9271_out0 = v_G1_8125_out0;
assign v_S_9273_out0 = v_G1_8127_out0;
assign v_S_9275_out0 = v_G1_8129_out0;
assign v_S_9278_out0 = v_G1_8132_out0;
assign v_S_9280_out0 = v_G1_8134_out0;
assign v_S_9282_out0 = v_G1_8136_out0;
assign v_S_9284_out0 = v_G1_8138_out0;
assign v_S_9286_out0 = v_G1_8140_out0;
assign v_S_9288_out0 = v_G1_8142_out0;
assign v_S_9290_out0 = v_G1_8144_out0;
assign v_S_9292_out0 = v_G1_8146_out0;
assign v_S_9294_out0 = v_G1_8148_out0;
assign v_S_9729_out0 = v_G1_8583_out0;
assign v_S_9731_out0 = v_G1_8585_out0;
assign v_S_9735_out0 = v_G1_8589_out0;
assign v_S_9737_out0 = v_G1_8591_out0;
assign v_S_9739_out0 = v_G1_8593_out0;
assign v_S_9742_out0 = v_G1_8596_out0;
assign v_S_9744_out0 = v_G1_8598_out0;
assign v_S_9746_out0 = v_G1_8600_out0;
assign v_S_9748_out0 = v_G1_8602_out0;
assign v_S_9750_out0 = v_G1_8604_out0;
assign v_S_9752_out0 = v_G1_8606_out0;
assign v_S_9754_out0 = v_G1_8608_out0;
assign v_S_9756_out0 = v_G1_8610_out0;
assign v_S_9758_out0 = v_G1_8612_out0;
assign v_CIN_10010_out0 = v_CARRY_5276_out0;
assign v_CIN_10234_out0 = v_CARRY_5740_out0;
assign v__681_out0 = { v__56_out0,v_S_4678_out0 };
assign v__682_out0 = { v__57_out0,v_S_4693_out0 };
assign v_RD_6282_out0 = v_CIN_10010_out0;
assign v_RD_6746_out0 = v_CIN_10234_out0;
assign v_RM_11705_out0 = v_S_9265_out0;
assign v_RM_11707_out0 = v_S_9267_out0;
assign v_RM_11711_out0 = v_S_9271_out0;
assign v_RM_11713_out0 = v_S_9273_out0;
assign v_RM_11715_out0 = v_S_9275_out0;
assign v_RM_11718_out0 = v_S_9278_out0;
assign v_RM_11720_out0 = v_S_9280_out0;
assign v_RM_11722_out0 = v_S_9282_out0;
assign v_RM_11724_out0 = v_S_9284_out0;
assign v_RM_11726_out0 = v_S_9286_out0;
assign v_RM_11728_out0 = v_S_9288_out0;
assign v_RM_11730_out0 = v_S_9290_out0;
assign v_RM_11732_out0 = v_S_9292_out0;
assign v_RM_11734_out0 = v_S_9294_out0;
assign v_RM_12169_out0 = v_S_9729_out0;
assign v_RM_12171_out0 = v_S_9731_out0;
assign v_RM_12175_out0 = v_S_9735_out0;
assign v_RM_12177_out0 = v_S_9737_out0;
assign v_RM_12179_out0 = v_S_9739_out0;
assign v_RM_12182_out0 = v_S_9742_out0;
assign v_RM_12184_out0 = v_S_9744_out0;
assign v_RM_12186_out0 = v_S_9746_out0;
assign v_RM_12188_out0 = v_S_9748_out0;
assign v_RM_12190_out0 = v_S_9750_out0;
assign v_RM_12192_out0 = v_S_9752_out0;
assign v_RM_12194_out0 = v_S_9754_out0;
assign v_RM_12196_out0 = v_S_9756_out0;
assign v_RM_12198_out0 = v_S_9758_out0;
assign v_G1_8137_out0 = ((v_RD_6282_out0 && !v_RM_11722_out0) || (!v_RD_6282_out0) && v_RM_11722_out0);
assign v_G1_8601_out0 = ((v_RD_6746_out0 && !v_RM_12186_out0) || (!v_RD_6746_out0) && v_RM_12186_out0);
assign v_G2_12673_out0 = v_RD_6282_out0 && v_RM_11722_out0;
assign v_G2_13137_out0 = v_RD_6746_out0 && v_RM_12186_out0;
assign v_CARRY_5282_out0 = v_G2_12673_out0;
assign v_CARRY_5746_out0 = v_G2_13137_out0;
assign v_S_9283_out0 = v_G1_8137_out0;
assign v_S_9747_out0 = v_G1_8601_out0;
assign v_S_1421_out0 = v_S_9283_out0;
assign v_S_1645_out0 = v_S_9747_out0;
assign v_G1_4197_out0 = v_CARRY_5282_out0 || v_CARRY_5281_out0;
assign v_G1_4421_out0 = v_CARRY_5746_out0 || v_CARRY_5745_out0;
assign v_COUT_889_out0 = v_G1_4197_out0;
assign v_COUT_1113_out0 = v_G1_4421_out0;
assign v_CIN_10016_out0 = v_COUT_889_out0;
assign v_CIN_10240_out0 = v_COUT_1113_out0;
assign v_RD_6294_out0 = v_CIN_10016_out0;
assign v_RD_6758_out0 = v_CIN_10240_out0;
assign v_G1_8149_out0 = ((v_RD_6294_out0 && !v_RM_11734_out0) || (!v_RD_6294_out0) && v_RM_11734_out0);
assign v_G1_8613_out0 = ((v_RD_6758_out0 && !v_RM_12198_out0) || (!v_RD_6758_out0) && v_RM_12198_out0);
assign v_G2_12685_out0 = v_RD_6294_out0 && v_RM_11734_out0;
assign v_G2_13149_out0 = v_RD_6758_out0 && v_RM_12198_out0;
assign v_CARRY_5294_out0 = v_G2_12685_out0;
assign v_CARRY_5758_out0 = v_G2_13149_out0;
assign v_S_9295_out0 = v_G1_8149_out0;
assign v_S_9759_out0 = v_G1_8613_out0;
assign v_S_1427_out0 = v_S_9295_out0;
assign v_S_1651_out0 = v_S_9759_out0;
assign v_G1_4203_out0 = v_CARRY_5294_out0 || v_CARRY_5293_out0;
assign v_G1_4427_out0 = v_CARRY_5758_out0 || v_CARRY_5757_out0;
assign v_COUT_895_out0 = v_G1_4203_out0;
assign v_COUT_1119_out0 = v_G1_4427_out0;
assign v__4795_out0 = { v_S_1421_out0,v_S_1427_out0 };
assign v__4810_out0 = { v_S_1645_out0,v_S_1651_out0 };
assign v_CIN_10011_out0 = v_COUT_895_out0;
assign v_CIN_10235_out0 = v_COUT_1119_out0;
assign v_RD_6284_out0 = v_CIN_10011_out0;
assign v_RD_6748_out0 = v_CIN_10235_out0;
assign v_G1_8139_out0 = ((v_RD_6284_out0 && !v_RM_11724_out0) || (!v_RD_6284_out0) && v_RM_11724_out0);
assign v_G1_8603_out0 = ((v_RD_6748_out0 && !v_RM_12188_out0) || (!v_RD_6748_out0) && v_RM_12188_out0);
assign v_G2_12675_out0 = v_RD_6284_out0 && v_RM_11724_out0;
assign v_G2_13139_out0 = v_RD_6748_out0 && v_RM_12188_out0;
assign v_CARRY_5284_out0 = v_G2_12675_out0;
assign v_CARRY_5748_out0 = v_G2_13139_out0;
assign v_S_9285_out0 = v_G1_8139_out0;
assign v_S_9749_out0 = v_G1_8603_out0;
assign v_S_1422_out0 = v_S_9285_out0;
assign v_S_1646_out0 = v_S_9749_out0;
assign v_G1_4198_out0 = v_CARRY_5284_out0 || v_CARRY_5283_out0;
assign v_G1_4422_out0 = v_CARRY_5748_out0 || v_CARRY_5747_out0;
assign v_COUT_890_out0 = v_G1_4198_out0;
assign v_COUT_1114_out0 = v_G1_4422_out0;
assign v__2565_out0 = { v__4795_out0,v_S_1422_out0 };
assign v__2580_out0 = { v__4810_out0,v_S_1646_out0 };
assign v_CIN_10006_out0 = v_COUT_890_out0;
assign v_CIN_10230_out0 = v_COUT_1114_out0;
assign v_RD_6273_out0 = v_CIN_10006_out0;
assign v_RD_6737_out0 = v_CIN_10230_out0;
assign v_G1_8128_out0 = ((v_RD_6273_out0 && !v_RM_11713_out0) || (!v_RD_6273_out0) && v_RM_11713_out0);
assign v_G1_8592_out0 = ((v_RD_6737_out0 && !v_RM_12177_out0) || (!v_RD_6737_out0) && v_RM_12177_out0);
assign v_G2_12664_out0 = v_RD_6273_out0 && v_RM_11713_out0;
assign v_G2_13128_out0 = v_RD_6737_out0 && v_RM_12177_out0;
assign v_CARRY_5273_out0 = v_G2_12664_out0;
assign v_CARRY_5737_out0 = v_G2_13128_out0;
assign v_S_9274_out0 = v_G1_8128_out0;
assign v_S_9738_out0 = v_G1_8592_out0;
assign v_S_1417_out0 = v_S_9274_out0;
assign v_S_1641_out0 = v_S_9738_out0;
assign v_G1_4193_out0 = v_CARRY_5273_out0 || v_CARRY_5272_out0;
assign v_G1_4417_out0 = v_CARRY_5737_out0 || v_CARRY_5736_out0;
assign v_COUT_885_out0 = v_G1_4193_out0;
assign v_COUT_1109_out0 = v_G1_4417_out0;
assign v__7045_out0 = { v__2565_out0,v_S_1417_out0 };
assign v__7060_out0 = { v__2580_out0,v_S_1641_out0 };
assign v_CIN_10005_out0 = v_COUT_885_out0;
assign v_CIN_10229_out0 = v_COUT_1109_out0;
assign v_RD_6271_out0 = v_CIN_10005_out0;
assign v_RD_6735_out0 = v_CIN_10229_out0;
assign v_G1_8126_out0 = ((v_RD_6271_out0 && !v_RM_11711_out0) || (!v_RD_6271_out0) && v_RM_11711_out0);
assign v_G1_8590_out0 = ((v_RD_6735_out0 && !v_RM_12175_out0) || (!v_RD_6735_out0) && v_RM_12175_out0);
assign v_G2_12662_out0 = v_RD_6271_out0 && v_RM_11711_out0;
assign v_G2_13126_out0 = v_RD_6735_out0 && v_RM_12175_out0;
assign v_CARRY_5271_out0 = v_G2_12662_out0;
assign v_CARRY_5735_out0 = v_G2_13126_out0;
assign v_S_9272_out0 = v_G1_8126_out0;
assign v_S_9736_out0 = v_G1_8590_out0;
assign v_S_1416_out0 = v_S_9272_out0;
assign v_S_1640_out0 = v_S_9736_out0;
assign v_G1_4192_out0 = v_CARRY_5271_out0 || v_CARRY_5270_out0;
assign v_G1_4416_out0 = v_CARRY_5735_out0 || v_CARRY_5734_out0;
assign v_COUT_884_out0 = v_G1_4192_out0;
assign v_COUT_1108_out0 = v_G1_4416_out0;
assign v__13531_out0 = { v__7045_out0,v_S_1416_out0 };
assign v__13546_out0 = { v__7060_out0,v_S_1640_out0 };
assign v_CIN_10012_out0 = v_COUT_884_out0;
assign v_CIN_10236_out0 = v_COUT_1108_out0;
assign v_RD_6286_out0 = v_CIN_10012_out0;
assign v_RD_6750_out0 = v_CIN_10236_out0;
assign v_G1_8141_out0 = ((v_RD_6286_out0 && !v_RM_11726_out0) || (!v_RD_6286_out0) && v_RM_11726_out0);
assign v_G1_8605_out0 = ((v_RD_6750_out0 && !v_RM_12190_out0) || (!v_RD_6750_out0) && v_RM_12190_out0);
assign v_G2_12677_out0 = v_RD_6286_out0 && v_RM_11726_out0;
assign v_G2_13141_out0 = v_RD_6750_out0 && v_RM_12190_out0;
assign v_CARRY_5286_out0 = v_G2_12677_out0;
assign v_CARRY_5750_out0 = v_G2_13141_out0;
assign v_S_9287_out0 = v_G1_8141_out0;
assign v_S_9751_out0 = v_G1_8605_out0;
assign v_S_1423_out0 = v_S_9287_out0;
assign v_S_1647_out0 = v_S_9751_out0;
assign v_G1_4199_out0 = v_CARRY_5286_out0 || v_CARRY_5285_out0;
assign v_G1_4423_out0 = v_CARRY_5750_out0 || v_CARRY_5749_out0;
assign v_COUT_891_out0 = v_G1_4199_out0;
assign v_COUT_1115_out0 = v_G1_4423_out0;
assign v__3324_out0 = { v__13531_out0,v_S_1423_out0 };
assign v__3339_out0 = { v__13546_out0,v_S_1647_out0 };
assign v_CIN_10013_out0 = v_COUT_891_out0;
assign v_CIN_10237_out0 = v_COUT_1115_out0;
assign v_RD_6288_out0 = v_CIN_10013_out0;
assign v_RD_6752_out0 = v_CIN_10237_out0;
assign v_G1_8143_out0 = ((v_RD_6288_out0 && !v_RM_11728_out0) || (!v_RD_6288_out0) && v_RM_11728_out0);
assign v_G1_8607_out0 = ((v_RD_6752_out0 && !v_RM_12192_out0) || (!v_RD_6752_out0) && v_RM_12192_out0);
assign v_G2_12679_out0 = v_RD_6288_out0 && v_RM_11728_out0;
assign v_G2_13143_out0 = v_RD_6752_out0 && v_RM_12192_out0;
assign v_CARRY_5288_out0 = v_G2_12679_out0;
assign v_CARRY_5752_out0 = v_G2_13143_out0;
assign v_S_9289_out0 = v_G1_8143_out0;
assign v_S_9753_out0 = v_G1_8607_out0;
assign v_S_1424_out0 = v_S_9289_out0;
assign v_S_1648_out0 = v_S_9753_out0;
assign v_G1_4200_out0 = v_CARRY_5288_out0 || v_CARRY_5287_out0;
assign v_G1_4424_out0 = v_CARRY_5752_out0 || v_CARRY_5751_out0;
assign v_COUT_892_out0 = v_G1_4200_out0;
assign v_COUT_1116_out0 = v_G1_4424_out0;
assign v__7160_out0 = { v__3324_out0,v_S_1424_out0 };
assign v__7175_out0 = { v__3339_out0,v_S_1648_out0 };
assign v_CIN_10015_out0 = v_COUT_892_out0;
assign v_CIN_10239_out0 = v_COUT_1116_out0;
assign v_RD_6292_out0 = v_CIN_10015_out0;
assign v_RD_6756_out0 = v_CIN_10239_out0;
assign v_G1_8147_out0 = ((v_RD_6292_out0 && !v_RM_11732_out0) || (!v_RD_6292_out0) && v_RM_11732_out0);
assign v_G1_8611_out0 = ((v_RD_6756_out0 && !v_RM_12196_out0) || (!v_RD_6756_out0) && v_RM_12196_out0);
assign v_G2_12683_out0 = v_RD_6292_out0 && v_RM_11732_out0;
assign v_G2_13147_out0 = v_RD_6756_out0 && v_RM_12196_out0;
assign v_CARRY_5292_out0 = v_G2_12683_out0;
assign v_CARRY_5756_out0 = v_G2_13147_out0;
assign v_S_9293_out0 = v_G1_8147_out0;
assign v_S_9757_out0 = v_G1_8611_out0;
assign v_S_1426_out0 = v_S_9293_out0;
assign v_S_1650_out0 = v_S_9757_out0;
assign v_G1_4202_out0 = v_CARRY_5292_out0 || v_CARRY_5291_out0;
assign v_G1_4426_out0 = v_CARRY_5756_out0 || v_CARRY_5755_out0;
assign v_COUT_894_out0 = v_G1_4202_out0;
assign v_COUT_1118_out0 = v_G1_4426_out0;
assign v__4762_out0 = { v__7160_out0,v_S_1426_out0 };
assign v__4777_out0 = { v__7175_out0,v_S_1650_out0 };
assign v_CIN_10008_out0 = v_COUT_894_out0;
assign v_CIN_10232_out0 = v_COUT_1118_out0;
assign v_RD_6278_out0 = v_CIN_10008_out0;
assign v_RD_6742_out0 = v_CIN_10232_out0;
assign v_G1_8133_out0 = ((v_RD_6278_out0 && !v_RM_11718_out0) || (!v_RD_6278_out0) && v_RM_11718_out0);
assign v_G1_8597_out0 = ((v_RD_6742_out0 && !v_RM_12182_out0) || (!v_RD_6742_out0) && v_RM_12182_out0);
assign v_G2_12669_out0 = v_RD_6278_out0 && v_RM_11718_out0;
assign v_G2_13133_out0 = v_RD_6742_out0 && v_RM_12182_out0;
assign v_CARRY_5278_out0 = v_G2_12669_out0;
assign v_CARRY_5742_out0 = v_G2_13133_out0;
assign v_S_9279_out0 = v_G1_8133_out0;
assign v_S_9743_out0 = v_G1_8597_out0;
assign v_S_1419_out0 = v_S_9279_out0;
assign v_S_1643_out0 = v_S_9743_out0;
assign v_G1_4195_out0 = v_CARRY_5278_out0 || v_CARRY_5277_out0;
assign v_G1_4419_out0 = v_CARRY_5742_out0 || v_CARRY_5741_out0;
assign v_COUT_887_out0 = v_G1_4195_out0;
assign v_COUT_1111_out0 = v_G1_4419_out0;
assign v__6939_out0 = { v__4762_out0,v_S_1419_out0 };
assign v__6954_out0 = { v__4777_out0,v_S_1643_out0 };
assign v_CIN_10009_out0 = v_COUT_887_out0;
assign v_CIN_10233_out0 = v_COUT_1111_out0;
assign v_RD_6280_out0 = v_CIN_10009_out0;
assign v_RD_6744_out0 = v_CIN_10233_out0;
assign v_G1_8135_out0 = ((v_RD_6280_out0 && !v_RM_11720_out0) || (!v_RD_6280_out0) && v_RM_11720_out0);
assign v_G1_8599_out0 = ((v_RD_6744_out0 && !v_RM_12184_out0) || (!v_RD_6744_out0) && v_RM_12184_out0);
assign v_G2_12671_out0 = v_RD_6280_out0 && v_RM_11720_out0;
assign v_G2_13135_out0 = v_RD_6744_out0 && v_RM_12184_out0;
assign v_CARRY_5280_out0 = v_G2_12671_out0;
assign v_CARRY_5744_out0 = v_G2_13135_out0;
assign v_S_9281_out0 = v_G1_8135_out0;
assign v_S_9745_out0 = v_G1_8599_out0;
assign v_S_1420_out0 = v_S_9281_out0;
assign v_S_1644_out0 = v_S_9745_out0;
assign v_G1_4196_out0 = v_CARRY_5280_out0 || v_CARRY_5279_out0;
assign v_G1_4420_out0 = v_CARRY_5744_out0 || v_CARRY_5743_out0;
assign v_COUT_888_out0 = v_G1_4196_out0;
assign v_COUT_1112_out0 = v_G1_4420_out0;
assign v__5815_out0 = { v__6939_out0,v_S_1420_out0 };
assign v__5830_out0 = { v__6954_out0,v_S_1644_out0 };
assign v_CIN_10014_out0 = v_COUT_888_out0;
assign v_CIN_10238_out0 = v_COUT_1112_out0;
assign v_RD_6290_out0 = v_CIN_10014_out0;
assign v_RD_6754_out0 = v_CIN_10238_out0;
assign v_G1_8145_out0 = ((v_RD_6290_out0 && !v_RM_11730_out0) || (!v_RD_6290_out0) && v_RM_11730_out0);
assign v_G1_8609_out0 = ((v_RD_6754_out0 && !v_RM_12194_out0) || (!v_RD_6754_out0) && v_RM_12194_out0);
assign v_G2_12681_out0 = v_RD_6290_out0 && v_RM_11730_out0;
assign v_G2_13145_out0 = v_RD_6754_out0 && v_RM_12194_out0;
assign v_CARRY_5290_out0 = v_G2_12681_out0;
assign v_CARRY_5754_out0 = v_G2_13145_out0;
assign v_S_9291_out0 = v_G1_8145_out0;
assign v_S_9755_out0 = v_G1_8609_out0;
assign v_S_1425_out0 = v_S_9291_out0;
assign v_S_1649_out0 = v_S_9755_out0;
assign v_G1_4201_out0 = v_CARRY_5290_out0 || v_CARRY_5289_out0;
assign v_G1_4425_out0 = v_CARRY_5754_out0 || v_CARRY_5753_out0;
assign v_COUT_893_out0 = v_G1_4201_out0;
assign v_COUT_1117_out0 = v_G1_4425_out0;
assign v__2039_out0 = { v__5815_out0,v_S_1425_out0 };
assign v__2054_out0 = { v__5830_out0,v_S_1649_out0 };
assign v_CIN_10002_out0 = v_COUT_893_out0;
assign v_CIN_10226_out0 = v_COUT_1117_out0;
assign v_RD_6265_out0 = v_CIN_10002_out0;
assign v_RD_6729_out0 = v_CIN_10226_out0;
assign v_G1_8120_out0 = ((v_RD_6265_out0 && !v_RM_11705_out0) || (!v_RD_6265_out0) && v_RM_11705_out0);
assign v_G1_8584_out0 = ((v_RD_6729_out0 && !v_RM_12169_out0) || (!v_RD_6729_out0) && v_RM_12169_out0);
assign v_G2_12656_out0 = v_RD_6265_out0 && v_RM_11705_out0;
assign v_G2_13120_out0 = v_RD_6729_out0 && v_RM_12169_out0;
assign v_CARRY_5265_out0 = v_G2_12656_out0;
assign v_CARRY_5729_out0 = v_G2_13120_out0;
assign v_S_9266_out0 = v_G1_8120_out0;
assign v_S_9730_out0 = v_G1_8584_out0;
assign v_S_1413_out0 = v_S_9266_out0;
assign v_S_1637_out0 = v_S_9730_out0;
assign v_G1_4189_out0 = v_CARRY_5265_out0 || v_CARRY_5264_out0;
assign v_G1_4413_out0 = v_CARRY_5729_out0 || v_CARRY_5728_out0;
assign v_COUT_881_out0 = v_G1_4189_out0;
assign v_COUT_1105_out0 = v_G1_4413_out0;
assign v__2806_out0 = { v__2039_out0,v_S_1413_out0 };
assign v__2821_out0 = { v__2054_out0,v_S_1637_out0 };
assign v_CIN_10007_out0 = v_COUT_881_out0;
assign v_CIN_10231_out0 = v_COUT_1105_out0;
assign v_RD_6275_out0 = v_CIN_10007_out0;
assign v_RD_6739_out0 = v_CIN_10231_out0;
assign v_G1_8130_out0 = ((v_RD_6275_out0 && !v_RM_11715_out0) || (!v_RD_6275_out0) && v_RM_11715_out0);
assign v_G1_8594_out0 = ((v_RD_6739_out0 && !v_RM_12179_out0) || (!v_RD_6739_out0) && v_RM_12179_out0);
assign v_G2_12666_out0 = v_RD_6275_out0 && v_RM_11715_out0;
assign v_G2_13130_out0 = v_RD_6739_out0 && v_RM_12179_out0;
assign v_CARRY_5275_out0 = v_G2_12666_out0;
assign v_CARRY_5739_out0 = v_G2_13130_out0;
assign v_S_9276_out0 = v_G1_8130_out0;
assign v_S_9740_out0 = v_G1_8594_out0;
assign v_S_1418_out0 = v_S_9276_out0;
assign v_S_1642_out0 = v_S_9740_out0;
assign v_G1_4194_out0 = v_CARRY_5275_out0 || v_CARRY_5274_out0;
assign v_G1_4418_out0 = v_CARRY_5739_out0 || v_CARRY_5738_out0;
assign v_COUT_886_out0 = v_G1_4194_out0;
assign v_COUT_1110_out0 = v_G1_4418_out0;
assign v__1838_out0 = { v__2806_out0,v_S_1418_out0 };
assign v__1853_out0 = { v__2821_out0,v_S_1642_out0 };
assign v_CIN_10003_out0 = v_COUT_886_out0;
assign v_CIN_10227_out0 = v_COUT_1110_out0;
assign v_RD_6267_out0 = v_CIN_10003_out0;
assign v_RD_6731_out0 = v_CIN_10227_out0;
assign v_G1_8122_out0 = ((v_RD_6267_out0 && !v_RM_11707_out0) || (!v_RD_6267_out0) && v_RM_11707_out0);
assign v_G1_8586_out0 = ((v_RD_6731_out0 && !v_RM_12171_out0) || (!v_RD_6731_out0) && v_RM_12171_out0);
assign v_G2_12658_out0 = v_RD_6267_out0 && v_RM_11707_out0;
assign v_G2_13122_out0 = v_RD_6731_out0 && v_RM_12171_out0;
assign v_CARRY_5267_out0 = v_G2_12658_out0;
assign v_CARRY_5731_out0 = v_G2_13122_out0;
assign v_S_9268_out0 = v_G1_8122_out0;
assign v_S_9732_out0 = v_G1_8586_out0;
assign v_S_1414_out0 = v_S_9268_out0;
assign v_S_1638_out0 = v_S_9732_out0;
assign v_G1_4190_out0 = v_CARRY_5267_out0 || v_CARRY_5266_out0;
assign v_G1_4414_out0 = v_CARRY_5731_out0 || v_CARRY_5730_out0;
assign v_COUT_882_out0 = v_G1_4190_out0;
assign v_COUT_1106_out0 = v_G1_4414_out0;
assign v__4562_out0 = { v__1838_out0,v_S_1414_out0 };
assign v__4577_out0 = { v__1853_out0,v_S_1638_out0 };
assign v_RM_3551_out0 = v_COUT_882_out0;
assign v_RM_3775_out0 = v_COUT_1106_out0;
assign v_RM_11708_out0 = v_RM_3551_out0;
assign v_RM_12172_out0 = v_RM_3775_out0;
assign v_G1_8123_out0 = ((v_RD_6268_out0 && !v_RM_11708_out0) || (!v_RD_6268_out0) && v_RM_11708_out0);
assign v_G1_8587_out0 = ((v_RD_6732_out0 && !v_RM_12172_out0) || (!v_RD_6732_out0) && v_RM_12172_out0);
assign v_G2_12659_out0 = v_RD_6268_out0 && v_RM_11708_out0;
assign v_G2_13123_out0 = v_RD_6732_out0 && v_RM_12172_out0;
assign v_CARRY_5268_out0 = v_G2_12659_out0;
assign v_CARRY_5732_out0 = v_G2_13123_out0;
assign v_S_9269_out0 = v_G1_8123_out0;
assign v_S_9733_out0 = v_G1_8587_out0;
assign v_RM_11709_out0 = v_S_9269_out0;
assign v_RM_12173_out0 = v_S_9733_out0;
assign v_G1_8124_out0 = ((v_RD_6269_out0 && !v_RM_11709_out0) || (!v_RD_6269_out0) && v_RM_11709_out0);
assign v_G1_8588_out0 = ((v_RD_6733_out0 && !v_RM_12173_out0) || (!v_RD_6733_out0) && v_RM_12173_out0);
assign v_G2_12660_out0 = v_RD_6269_out0 && v_RM_11709_out0;
assign v_G2_13124_out0 = v_RD_6733_out0 && v_RM_12173_out0;
assign v_CARRY_5269_out0 = v_G2_12660_out0;
assign v_CARRY_5733_out0 = v_G2_13124_out0;
assign v_S_9270_out0 = v_G1_8124_out0;
assign v_S_9734_out0 = v_G1_8588_out0;
assign v_S_1415_out0 = v_S_9270_out0;
assign v_S_1639_out0 = v_S_9734_out0;
assign v_G1_4191_out0 = v_CARRY_5269_out0 || v_CARRY_5268_out0;
assign v_G1_4415_out0 = v_CARRY_5733_out0 || v_CARRY_5732_out0;
assign v_COUT_883_out0 = v_G1_4191_out0;
assign v_COUT_1107_out0 = v_G1_4415_out0;
assign v__10664_out0 = { v__4562_out0,v_S_1415_out0 };
assign v__10679_out0 = { v__4577_out0,v_S_1639_out0 };
assign v__10959_out0 = { v__10664_out0,v_COUT_883_out0 };
assign v__10974_out0 = { v__10679_out0,v_COUT_1107_out0 };
assign v_COUT_10929_out0 = v__10959_out0;
assign v_COUT_10944_out0 = v__10974_out0;
assign v_CIN_2366_out0 = v_COUT_10929_out0;
assign v_CIN_2381_out0 = v_COUT_10944_out0;
assign v__479_out0 = v_CIN_2366_out0[8:8];
assign v__494_out0 = v_CIN_2381_out0[8:8];
assign v__1784_out0 = v_CIN_2366_out0[6:6];
assign v__1799_out0 = v_CIN_2381_out0[6:6];
assign v__2166_out0 = v_CIN_2366_out0[3:3];
assign v__2181_out0 = v_CIN_2381_out0[3:3];
assign v__2205_out0 = v_CIN_2366_out0[15:15];
assign v__2219_out0 = v_CIN_2381_out0[15:15];
assign v__2513_out0 = v_CIN_2366_out0[0:0];
assign v__2528_out0 = v_CIN_2381_out0[0:0];
assign v__3062_out0 = v_CIN_2366_out0[9:9];
assign v__3077_out0 = v_CIN_2381_out0[9:9];
assign v__3096_out0 = v_CIN_2366_out0[2:2];
assign v__3111_out0 = v_CIN_2381_out0[2:2];
assign v__3150_out0 = v_CIN_2366_out0[7:7];
assign v__3165_out0 = v_CIN_2381_out0[7:7];
assign v__3834_out0 = v_CIN_2366_out0[1:1];
assign v__3849_out0 = v_CIN_2381_out0[1:1];
assign v__3872_out0 = v_CIN_2366_out0[10:10];
assign v__3887_out0 = v_CIN_2381_out0[10:10];
assign v__6811_out0 = v_CIN_2366_out0[11:11];
assign v__6826_out0 = v_CIN_2381_out0[11:11];
assign v__7655_out0 = v_CIN_2366_out0[12:12];
assign v__7670_out0 = v_CIN_2381_out0[12:12];
assign v__8710_out0 = v_CIN_2366_out0[13:13];
assign v__8725_out0 = v_CIN_2381_out0[13:13];
assign v__8780_out0 = v_CIN_2366_out0[14:14];
assign v__8795_out0 = v_CIN_2381_out0[14:14];
assign v__10730_out0 = v_CIN_2366_out0[5:5];
assign v__10745_out0 = v_CIN_2381_out0[5:5];
assign v__13459_out0 = v_CIN_2366_out0[4:4];
assign v__13474_out0 = v_CIN_2381_out0[4:4];
assign v_RM_3519_out0 = v__7655_out0;
assign v_RM_3520_out0 = v__8780_out0;
assign v_RM_3522_out0 = v__10730_out0;
assign v_RM_3523_out0 = v__13459_out0;
assign v_RM_3524_out0 = v__8710_out0;
assign v_RM_3525_out0 = v__3062_out0;
assign v_RM_3526_out0 = v__3872_out0;
assign v_RM_3527_out0 = v__3834_out0;
assign v_RM_3528_out0 = v__2166_out0;
assign v_RM_3529_out0 = v__1784_out0;
assign v_RM_3530_out0 = v__3150_out0;
assign v_RM_3531_out0 = v__6811_out0;
assign v_RM_3532_out0 = v__479_out0;
assign v_RM_3533_out0 = v__3096_out0;
assign v_RM_3743_out0 = v__7670_out0;
assign v_RM_3744_out0 = v__8795_out0;
assign v_RM_3746_out0 = v__10745_out0;
assign v_RM_3747_out0 = v__13474_out0;
assign v_RM_3748_out0 = v__8725_out0;
assign v_RM_3749_out0 = v__3077_out0;
assign v_RM_3750_out0 = v__3887_out0;
assign v_RM_3751_out0 = v__3849_out0;
assign v_RM_3752_out0 = v__2181_out0;
assign v_RM_3753_out0 = v__1799_out0;
assign v_RM_3754_out0 = v__3165_out0;
assign v_RM_3755_out0 = v__6826_out0;
assign v_RM_3756_out0 = v__494_out0;
assign v_RM_3757_out0 = v__3111_out0;
assign v_CIN_9974_out0 = v__2205_out0;
assign v_CIN_10198_out0 = v__2219_out0;
assign v_RM_11654_out0 = v__2513_out0;
assign v_RM_12118_out0 = v__2528_out0;
assign v_RD_6207_out0 = v_CIN_9974_out0;
assign v_RD_6671_out0 = v_CIN_10198_out0;
assign v_G1_8069_out0 = ((v_RD_6214_out0 && !v_RM_11654_out0) || (!v_RD_6214_out0) && v_RM_11654_out0);
assign v_G1_8533_out0 = ((v_RD_6678_out0 && !v_RM_12118_out0) || (!v_RD_6678_out0) && v_RM_12118_out0);
assign v_RM_11642_out0 = v_RM_3519_out0;
assign v_RM_11644_out0 = v_RM_3520_out0;
assign v_RM_11648_out0 = v_RM_3522_out0;
assign v_RM_11650_out0 = v_RM_3523_out0;
assign v_RM_11652_out0 = v_RM_3524_out0;
assign v_RM_11655_out0 = v_RM_3525_out0;
assign v_RM_11657_out0 = v_RM_3526_out0;
assign v_RM_11659_out0 = v_RM_3527_out0;
assign v_RM_11661_out0 = v_RM_3528_out0;
assign v_RM_11663_out0 = v_RM_3529_out0;
assign v_RM_11665_out0 = v_RM_3530_out0;
assign v_RM_11667_out0 = v_RM_3531_out0;
assign v_RM_11669_out0 = v_RM_3532_out0;
assign v_RM_11671_out0 = v_RM_3533_out0;
assign v_RM_12106_out0 = v_RM_3743_out0;
assign v_RM_12108_out0 = v_RM_3744_out0;
assign v_RM_12112_out0 = v_RM_3746_out0;
assign v_RM_12114_out0 = v_RM_3747_out0;
assign v_RM_12116_out0 = v_RM_3748_out0;
assign v_RM_12119_out0 = v_RM_3749_out0;
assign v_RM_12121_out0 = v_RM_3750_out0;
assign v_RM_12123_out0 = v_RM_3751_out0;
assign v_RM_12125_out0 = v_RM_3752_out0;
assign v_RM_12127_out0 = v_RM_3753_out0;
assign v_RM_12129_out0 = v_RM_3754_out0;
assign v_RM_12131_out0 = v_RM_3755_out0;
assign v_RM_12133_out0 = v_RM_3756_out0;
assign v_RM_12135_out0 = v_RM_3757_out0;
assign v_G2_12605_out0 = v_RD_6214_out0 && v_RM_11654_out0;
assign v_G2_13069_out0 = v_RD_6678_out0 && v_RM_12118_out0;
assign v_CARRY_5214_out0 = v_G2_12605_out0;
assign v_CARRY_5678_out0 = v_G2_13069_out0;
assign v_G1_8057_out0 = ((v_RD_6202_out0 && !v_RM_11642_out0) || (!v_RD_6202_out0) && v_RM_11642_out0);
assign v_G1_8059_out0 = ((v_RD_6204_out0 && !v_RM_11644_out0) || (!v_RD_6204_out0) && v_RM_11644_out0);
assign v_G1_8063_out0 = ((v_RD_6208_out0 && !v_RM_11648_out0) || (!v_RD_6208_out0) && v_RM_11648_out0);
assign v_G1_8065_out0 = ((v_RD_6210_out0 && !v_RM_11650_out0) || (!v_RD_6210_out0) && v_RM_11650_out0);
assign v_G1_8067_out0 = ((v_RD_6212_out0 && !v_RM_11652_out0) || (!v_RD_6212_out0) && v_RM_11652_out0);
assign v_G1_8070_out0 = ((v_RD_6215_out0 && !v_RM_11655_out0) || (!v_RD_6215_out0) && v_RM_11655_out0);
assign v_G1_8072_out0 = ((v_RD_6217_out0 && !v_RM_11657_out0) || (!v_RD_6217_out0) && v_RM_11657_out0);
assign v_G1_8074_out0 = ((v_RD_6219_out0 && !v_RM_11659_out0) || (!v_RD_6219_out0) && v_RM_11659_out0);
assign v_G1_8076_out0 = ((v_RD_6221_out0 && !v_RM_11661_out0) || (!v_RD_6221_out0) && v_RM_11661_out0);
assign v_G1_8078_out0 = ((v_RD_6223_out0 && !v_RM_11663_out0) || (!v_RD_6223_out0) && v_RM_11663_out0);
assign v_G1_8080_out0 = ((v_RD_6225_out0 && !v_RM_11665_out0) || (!v_RD_6225_out0) && v_RM_11665_out0);
assign v_G1_8082_out0 = ((v_RD_6227_out0 && !v_RM_11667_out0) || (!v_RD_6227_out0) && v_RM_11667_out0);
assign v_G1_8084_out0 = ((v_RD_6229_out0 && !v_RM_11669_out0) || (!v_RD_6229_out0) && v_RM_11669_out0);
assign v_G1_8086_out0 = ((v_RD_6231_out0 && !v_RM_11671_out0) || (!v_RD_6231_out0) && v_RM_11671_out0);
assign v_G1_8521_out0 = ((v_RD_6666_out0 && !v_RM_12106_out0) || (!v_RD_6666_out0) && v_RM_12106_out0);
assign v_G1_8523_out0 = ((v_RD_6668_out0 && !v_RM_12108_out0) || (!v_RD_6668_out0) && v_RM_12108_out0);
assign v_G1_8527_out0 = ((v_RD_6672_out0 && !v_RM_12112_out0) || (!v_RD_6672_out0) && v_RM_12112_out0);
assign v_G1_8529_out0 = ((v_RD_6674_out0 && !v_RM_12114_out0) || (!v_RD_6674_out0) && v_RM_12114_out0);
assign v_G1_8531_out0 = ((v_RD_6676_out0 && !v_RM_12116_out0) || (!v_RD_6676_out0) && v_RM_12116_out0);
assign v_G1_8534_out0 = ((v_RD_6679_out0 && !v_RM_12119_out0) || (!v_RD_6679_out0) && v_RM_12119_out0);
assign v_G1_8536_out0 = ((v_RD_6681_out0 && !v_RM_12121_out0) || (!v_RD_6681_out0) && v_RM_12121_out0);
assign v_G1_8538_out0 = ((v_RD_6683_out0 && !v_RM_12123_out0) || (!v_RD_6683_out0) && v_RM_12123_out0);
assign v_G1_8540_out0 = ((v_RD_6685_out0 && !v_RM_12125_out0) || (!v_RD_6685_out0) && v_RM_12125_out0);
assign v_G1_8542_out0 = ((v_RD_6687_out0 && !v_RM_12127_out0) || (!v_RD_6687_out0) && v_RM_12127_out0);
assign v_G1_8544_out0 = ((v_RD_6689_out0 && !v_RM_12129_out0) || (!v_RD_6689_out0) && v_RM_12129_out0);
assign v_G1_8546_out0 = ((v_RD_6691_out0 && !v_RM_12131_out0) || (!v_RD_6691_out0) && v_RM_12131_out0);
assign v_G1_8548_out0 = ((v_RD_6693_out0 && !v_RM_12133_out0) || (!v_RD_6693_out0) && v_RM_12133_out0);
assign v_G1_8550_out0 = ((v_RD_6695_out0 && !v_RM_12135_out0) || (!v_RD_6695_out0) && v_RM_12135_out0);
assign v_S_9215_out0 = v_G1_8069_out0;
assign v_S_9679_out0 = v_G1_8533_out0;
assign v_G2_12593_out0 = v_RD_6202_out0 && v_RM_11642_out0;
assign v_G2_12595_out0 = v_RD_6204_out0 && v_RM_11644_out0;
assign v_G2_12599_out0 = v_RD_6208_out0 && v_RM_11648_out0;
assign v_G2_12601_out0 = v_RD_6210_out0 && v_RM_11650_out0;
assign v_G2_12603_out0 = v_RD_6212_out0 && v_RM_11652_out0;
assign v_G2_12606_out0 = v_RD_6215_out0 && v_RM_11655_out0;
assign v_G2_12608_out0 = v_RD_6217_out0 && v_RM_11657_out0;
assign v_G2_12610_out0 = v_RD_6219_out0 && v_RM_11659_out0;
assign v_G2_12612_out0 = v_RD_6221_out0 && v_RM_11661_out0;
assign v_G2_12614_out0 = v_RD_6223_out0 && v_RM_11663_out0;
assign v_G2_12616_out0 = v_RD_6225_out0 && v_RM_11665_out0;
assign v_G2_12618_out0 = v_RD_6227_out0 && v_RM_11667_out0;
assign v_G2_12620_out0 = v_RD_6229_out0 && v_RM_11669_out0;
assign v_G2_12622_out0 = v_RD_6231_out0 && v_RM_11671_out0;
assign v_G2_13057_out0 = v_RD_6666_out0 && v_RM_12106_out0;
assign v_G2_13059_out0 = v_RD_6668_out0 && v_RM_12108_out0;
assign v_G2_13063_out0 = v_RD_6672_out0 && v_RM_12112_out0;
assign v_G2_13065_out0 = v_RD_6674_out0 && v_RM_12114_out0;
assign v_G2_13067_out0 = v_RD_6676_out0 && v_RM_12116_out0;
assign v_G2_13070_out0 = v_RD_6679_out0 && v_RM_12119_out0;
assign v_G2_13072_out0 = v_RD_6681_out0 && v_RM_12121_out0;
assign v_G2_13074_out0 = v_RD_6683_out0 && v_RM_12123_out0;
assign v_G2_13076_out0 = v_RD_6685_out0 && v_RM_12125_out0;
assign v_G2_13078_out0 = v_RD_6687_out0 && v_RM_12127_out0;
assign v_G2_13080_out0 = v_RD_6689_out0 && v_RM_12129_out0;
assign v_G2_13082_out0 = v_RD_6691_out0 && v_RM_12131_out0;
assign v_G2_13084_out0 = v_RD_6693_out0 && v_RM_12133_out0;
assign v_G2_13086_out0 = v_RD_6695_out0 && v_RM_12135_out0;
assign v_S_4676_out0 = v_S_9215_out0;
assign v_S_4691_out0 = v_S_9679_out0;
assign v_CARRY_5202_out0 = v_G2_12593_out0;
assign v_CARRY_5204_out0 = v_G2_12595_out0;
assign v_CARRY_5208_out0 = v_G2_12599_out0;
assign v_CARRY_5210_out0 = v_G2_12601_out0;
assign v_CARRY_5212_out0 = v_G2_12603_out0;
assign v_CARRY_5215_out0 = v_G2_12606_out0;
assign v_CARRY_5217_out0 = v_G2_12608_out0;
assign v_CARRY_5219_out0 = v_G2_12610_out0;
assign v_CARRY_5221_out0 = v_G2_12612_out0;
assign v_CARRY_5223_out0 = v_G2_12614_out0;
assign v_CARRY_5225_out0 = v_G2_12616_out0;
assign v_CARRY_5227_out0 = v_G2_12618_out0;
assign v_CARRY_5229_out0 = v_G2_12620_out0;
assign v_CARRY_5231_out0 = v_G2_12622_out0;
assign v_CARRY_5666_out0 = v_G2_13057_out0;
assign v_CARRY_5668_out0 = v_G2_13059_out0;
assign v_CARRY_5672_out0 = v_G2_13063_out0;
assign v_CARRY_5674_out0 = v_G2_13065_out0;
assign v_CARRY_5676_out0 = v_G2_13067_out0;
assign v_CARRY_5679_out0 = v_G2_13070_out0;
assign v_CARRY_5681_out0 = v_G2_13072_out0;
assign v_CARRY_5683_out0 = v_G2_13074_out0;
assign v_CARRY_5685_out0 = v_G2_13076_out0;
assign v_CARRY_5687_out0 = v_G2_13078_out0;
assign v_CARRY_5689_out0 = v_G2_13080_out0;
assign v_CARRY_5691_out0 = v_G2_13082_out0;
assign v_CARRY_5693_out0 = v_G2_13084_out0;
assign v_CARRY_5695_out0 = v_G2_13086_out0;
assign v_S_9203_out0 = v_G1_8057_out0;
assign v_S_9205_out0 = v_G1_8059_out0;
assign v_S_9209_out0 = v_G1_8063_out0;
assign v_S_9211_out0 = v_G1_8065_out0;
assign v_S_9213_out0 = v_G1_8067_out0;
assign v_S_9216_out0 = v_G1_8070_out0;
assign v_S_9218_out0 = v_G1_8072_out0;
assign v_S_9220_out0 = v_G1_8074_out0;
assign v_S_9222_out0 = v_G1_8076_out0;
assign v_S_9224_out0 = v_G1_8078_out0;
assign v_S_9226_out0 = v_G1_8080_out0;
assign v_S_9228_out0 = v_G1_8082_out0;
assign v_S_9230_out0 = v_G1_8084_out0;
assign v_S_9232_out0 = v_G1_8086_out0;
assign v_S_9667_out0 = v_G1_8521_out0;
assign v_S_9669_out0 = v_G1_8523_out0;
assign v_S_9673_out0 = v_G1_8527_out0;
assign v_S_9675_out0 = v_G1_8529_out0;
assign v_S_9677_out0 = v_G1_8531_out0;
assign v_S_9680_out0 = v_G1_8534_out0;
assign v_S_9682_out0 = v_G1_8536_out0;
assign v_S_9684_out0 = v_G1_8538_out0;
assign v_S_9686_out0 = v_G1_8540_out0;
assign v_S_9688_out0 = v_G1_8542_out0;
assign v_S_9690_out0 = v_G1_8544_out0;
assign v_S_9692_out0 = v_G1_8546_out0;
assign v_S_9694_out0 = v_G1_8548_out0;
assign v_S_9696_out0 = v_G1_8550_out0;
assign v_CIN_9980_out0 = v_CARRY_5214_out0;
assign v_CIN_10204_out0 = v_CARRY_5678_out0;
assign v__636_out0 = { v__681_out0,v_S_4676_out0 };
assign v__637_out0 = { v__682_out0,v_S_4691_out0 };
assign v_RD_6220_out0 = v_CIN_9980_out0;
assign v_RD_6684_out0 = v_CIN_10204_out0;
assign v_RM_11643_out0 = v_S_9203_out0;
assign v_RM_11645_out0 = v_S_9205_out0;
assign v_RM_11649_out0 = v_S_9209_out0;
assign v_RM_11651_out0 = v_S_9211_out0;
assign v_RM_11653_out0 = v_S_9213_out0;
assign v_RM_11656_out0 = v_S_9216_out0;
assign v_RM_11658_out0 = v_S_9218_out0;
assign v_RM_11660_out0 = v_S_9220_out0;
assign v_RM_11662_out0 = v_S_9222_out0;
assign v_RM_11664_out0 = v_S_9224_out0;
assign v_RM_11666_out0 = v_S_9226_out0;
assign v_RM_11668_out0 = v_S_9228_out0;
assign v_RM_11670_out0 = v_S_9230_out0;
assign v_RM_11672_out0 = v_S_9232_out0;
assign v_RM_12107_out0 = v_S_9667_out0;
assign v_RM_12109_out0 = v_S_9669_out0;
assign v_RM_12113_out0 = v_S_9673_out0;
assign v_RM_12115_out0 = v_S_9675_out0;
assign v_RM_12117_out0 = v_S_9677_out0;
assign v_RM_12120_out0 = v_S_9680_out0;
assign v_RM_12122_out0 = v_S_9682_out0;
assign v_RM_12124_out0 = v_S_9684_out0;
assign v_RM_12126_out0 = v_S_9686_out0;
assign v_RM_12128_out0 = v_S_9688_out0;
assign v_RM_12130_out0 = v_S_9690_out0;
assign v_RM_12132_out0 = v_S_9692_out0;
assign v_RM_12134_out0 = v_S_9694_out0;
assign v_RM_12136_out0 = v_S_9696_out0;
assign v_G1_8075_out0 = ((v_RD_6220_out0 && !v_RM_11660_out0) || (!v_RD_6220_out0) && v_RM_11660_out0);
assign v_G1_8539_out0 = ((v_RD_6684_out0 && !v_RM_12124_out0) || (!v_RD_6684_out0) && v_RM_12124_out0);
assign v_G2_12611_out0 = v_RD_6220_out0 && v_RM_11660_out0;
assign v_G2_13075_out0 = v_RD_6684_out0 && v_RM_12124_out0;
assign v_CARRY_5220_out0 = v_G2_12611_out0;
assign v_CARRY_5684_out0 = v_G2_13075_out0;
assign v_S_9221_out0 = v_G1_8075_out0;
assign v_S_9685_out0 = v_G1_8539_out0;
assign v_S_1391_out0 = v_S_9221_out0;
assign v_S_1615_out0 = v_S_9685_out0;
assign v_G1_4167_out0 = v_CARRY_5220_out0 || v_CARRY_5219_out0;
assign v_G1_4391_out0 = v_CARRY_5684_out0 || v_CARRY_5683_out0;
assign v_COUT_859_out0 = v_G1_4167_out0;
assign v_COUT_1083_out0 = v_G1_4391_out0;
assign v_CIN_9986_out0 = v_COUT_859_out0;
assign v_CIN_10210_out0 = v_COUT_1083_out0;
assign v_RD_6232_out0 = v_CIN_9986_out0;
assign v_RD_6696_out0 = v_CIN_10210_out0;
assign v_G1_8087_out0 = ((v_RD_6232_out0 && !v_RM_11672_out0) || (!v_RD_6232_out0) && v_RM_11672_out0);
assign v_G1_8551_out0 = ((v_RD_6696_out0 && !v_RM_12136_out0) || (!v_RD_6696_out0) && v_RM_12136_out0);
assign v_G2_12623_out0 = v_RD_6232_out0 && v_RM_11672_out0;
assign v_G2_13087_out0 = v_RD_6696_out0 && v_RM_12136_out0;
assign v_CARRY_5232_out0 = v_G2_12623_out0;
assign v_CARRY_5696_out0 = v_G2_13087_out0;
assign v_S_9233_out0 = v_G1_8087_out0;
assign v_S_9697_out0 = v_G1_8551_out0;
assign v_S_1397_out0 = v_S_9233_out0;
assign v_S_1621_out0 = v_S_9697_out0;
assign v_G1_4173_out0 = v_CARRY_5232_out0 || v_CARRY_5231_out0;
assign v_G1_4397_out0 = v_CARRY_5696_out0 || v_CARRY_5695_out0;
assign v_COUT_865_out0 = v_G1_4173_out0;
assign v_COUT_1089_out0 = v_G1_4397_out0;
assign v__4793_out0 = { v_S_1391_out0,v_S_1397_out0 };
assign v__4808_out0 = { v_S_1615_out0,v_S_1621_out0 };
assign v_CIN_9981_out0 = v_COUT_865_out0;
assign v_CIN_10205_out0 = v_COUT_1089_out0;
assign v_RD_6222_out0 = v_CIN_9981_out0;
assign v_RD_6686_out0 = v_CIN_10205_out0;
assign v_G1_8077_out0 = ((v_RD_6222_out0 && !v_RM_11662_out0) || (!v_RD_6222_out0) && v_RM_11662_out0);
assign v_G1_8541_out0 = ((v_RD_6686_out0 && !v_RM_12126_out0) || (!v_RD_6686_out0) && v_RM_12126_out0);
assign v_G2_12613_out0 = v_RD_6222_out0 && v_RM_11662_out0;
assign v_G2_13077_out0 = v_RD_6686_out0 && v_RM_12126_out0;
assign v_CARRY_5222_out0 = v_G2_12613_out0;
assign v_CARRY_5686_out0 = v_G2_13077_out0;
assign v_S_9223_out0 = v_G1_8077_out0;
assign v_S_9687_out0 = v_G1_8541_out0;
assign v_S_1392_out0 = v_S_9223_out0;
assign v_S_1616_out0 = v_S_9687_out0;
assign v_G1_4168_out0 = v_CARRY_5222_out0 || v_CARRY_5221_out0;
assign v_G1_4392_out0 = v_CARRY_5686_out0 || v_CARRY_5685_out0;
assign v_COUT_860_out0 = v_G1_4168_out0;
assign v_COUT_1084_out0 = v_G1_4392_out0;
assign v__2563_out0 = { v__4793_out0,v_S_1392_out0 };
assign v__2578_out0 = { v__4808_out0,v_S_1616_out0 };
assign v_CIN_9976_out0 = v_COUT_860_out0;
assign v_CIN_10200_out0 = v_COUT_1084_out0;
assign v_RD_6211_out0 = v_CIN_9976_out0;
assign v_RD_6675_out0 = v_CIN_10200_out0;
assign v_G1_8066_out0 = ((v_RD_6211_out0 && !v_RM_11651_out0) || (!v_RD_6211_out0) && v_RM_11651_out0);
assign v_G1_8530_out0 = ((v_RD_6675_out0 && !v_RM_12115_out0) || (!v_RD_6675_out0) && v_RM_12115_out0);
assign v_G2_12602_out0 = v_RD_6211_out0 && v_RM_11651_out0;
assign v_G2_13066_out0 = v_RD_6675_out0 && v_RM_12115_out0;
assign v_CARRY_5211_out0 = v_G2_12602_out0;
assign v_CARRY_5675_out0 = v_G2_13066_out0;
assign v_S_9212_out0 = v_G1_8066_out0;
assign v_S_9676_out0 = v_G1_8530_out0;
assign v_S_1387_out0 = v_S_9212_out0;
assign v_S_1611_out0 = v_S_9676_out0;
assign v_G1_4163_out0 = v_CARRY_5211_out0 || v_CARRY_5210_out0;
assign v_G1_4387_out0 = v_CARRY_5675_out0 || v_CARRY_5674_out0;
assign v_COUT_855_out0 = v_G1_4163_out0;
assign v_COUT_1079_out0 = v_G1_4387_out0;
assign v__7043_out0 = { v__2563_out0,v_S_1387_out0 };
assign v__7058_out0 = { v__2578_out0,v_S_1611_out0 };
assign v_CIN_9975_out0 = v_COUT_855_out0;
assign v_CIN_10199_out0 = v_COUT_1079_out0;
assign v_RD_6209_out0 = v_CIN_9975_out0;
assign v_RD_6673_out0 = v_CIN_10199_out0;
assign v_G1_8064_out0 = ((v_RD_6209_out0 && !v_RM_11649_out0) || (!v_RD_6209_out0) && v_RM_11649_out0);
assign v_G1_8528_out0 = ((v_RD_6673_out0 && !v_RM_12113_out0) || (!v_RD_6673_out0) && v_RM_12113_out0);
assign v_G2_12600_out0 = v_RD_6209_out0 && v_RM_11649_out0;
assign v_G2_13064_out0 = v_RD_6673_out0 && v_RM_12113_out0;
assign v_CARRY_5209_out0 = v_G2_12600_out0;
assign v_CARRY_5673_out0 = v_G2_13064_out0;
assign v_S_9210_out0 = v_G1_8064_out0;
assign v_S_9674_out0 = v_G1_8528_out0;
assign v_S_1386_out0 = v_S_9210_out0;
assign v_S_1610_out0 = v_S_9674_out0;
assign v_G1_4162_out0 = v_CARRY_5209_out0 || v_CARRY_5208_out0;
assign v_G1_4386_out0 = v_CARRY_5673_out0 || v_CARRY_5672_out0;
assign v_COUT_854_out0 = v_G1_4162_out0;
assign v_COUT_1078_out0 = v_G1_4386_out0;
assign v__13529_out0 = { v__7043_out0,v_S_1386_out0 };
assign v__13544_out0 = { v__7058_out0,v_S_1610_out0 };
assign v_CIN_9982_out0 = v_COUT_854_out0;
assign v_CIN_10206_out0 = v_COUT_1078_out0;
assign v_RD_6224_out0 = v_CIN_9982_out0;
assign v_RD_6688_out0 = v_CIN_10206_out0;
assign v_G1_8079_out0 = ((v_RD_6224_out0 && !v_RM_11664_out0) || (!v_RD_6224_out0) && v_RM_11664_out0);
assign v_G1_8543_out0 = ((v_RD_6688_out0 && !v_RM_12128_out0) || (!v_RD_6688_out0) && v_RM_12128_out0);
assign v_G2_12615_out0 = v_RD_6224_out0 && v_RM_11664_out0;
assign v_G2_13079_out0 = v_RD_6688_out0 && v_RM_12128_out0;
assign v_CARRY_5224_out0 = v_G2_12615_out0;
assign v_CARRY_5688_out0 = v_G2_13079_out0;
assign v_S_9225_out0 = v_G1_8079_out0;
assign v_S_9689_out0 = v_G1_8543_out0;
assign v_S_1393_out0 = v_S_9225_out0;
assign v_S_1617_out0 = v_S_9689_out0;
assign v_G1_4169_out0 = v_CARRY_5224_out0 || v_CARRY_5223_out0;
assign v_G1_4393_out0 = v_CARRY_5688_out0 || v_CARRY_5687_out0;
assign v_COUT_861_out0 = v_G1_4169_out0;
assign v_COUT_1085_out0 = v_G1_4393_out0;
assign v__3322_out0 = { v__13529_out0,v_S_1393_out0 };
assign v__3337_out0 = { v__13544_out0,v_S_1617_out0 };
assign v_CIN_9983_out0 = v_COUT_861_out0;
assign v_CIN_10207_out0 = v_COUT_1085_out0;
assign v_RD_6226_out0 = v_CIN_9983_out0;
assign v_RD_6690_out0 = v_CIN_10207_out0;
assign v_G1_8081_out0 = ((v_RD_6226_out0 && !v_RM_11666_out0) || (!v_RD_6226_out0) && v_RM_11666_out0);
assign v_G1_8545_out0 = ((v_RD_6690_out0 && !v_RM_12130_out0) || (!v_RD_6690_out0) && v_RM_12130_out0);
assign v_G2_12617_out0 = v_RD_6226_out0 && v_RM_11666_out0;
assign v_G2_13081_out0 = v_RD_6690_out0 && v_RM_12130_out0;
assign v_CARRY_5226_out0 = v_G2_12617_out0;
assign v_CARRY_5690_out0 = v_G2_13081_out0;
assign v_S_9227_out0 = v_G1_8081_out0;
assign v_S_9691_out0 = v_G1_8545_out0;
assign v_S_1394_out0 = v_S_9227_out0;
assign v_S_1618_out0 = v_S_9691_out0;
assign v_G1_4170_out0 = v_CARRY_5226_out0 || v_CARRY_5225_out0;
assign v_G1_4394_out0 = v_CARRY_5690_out0 || v_CARRY_5689_out0;
assign v_COUT_862_out0 = v_G1_4170_out0;
assign v_COUT_1086_out0 = v_G1_4394_out0;
assign v__7158_out0 = { v__3322_out0,v_S_1394_out0 };
assign v__7173_out0 = { v__3337_out0,v_S_1618_out0 };
assign v_CIN_9985_out0 = v_COUT_862_out0;
assign v_CIN_10209_out0 = v_COUT_1086_out0;
assign v_RD_6230_out0 = v_CIN_9985_out0;
assign v_RD_6694_out0 = v_CIN_10209_out0;
assign v_G1_8085_out0 = ((v_RD_6230_out0 && !v_RM_11670_out0) || (!v_RD_6230_out0) && v_RM_11670_out0);
assign v_G1_8549_out0 = ((v_RD_6694_out0 && !v_RM_12134_out0) || (!v_RD_6694_out0) && v_RM_12134_out0);
assign v_G2_12621_out0 = v_RD_6230_out0 && v_RM_11670_out0;
assign v_G2_13085_out0 = v_RD_6694_out0 && v_RM_12134_out0;
assign v_CARRY_5230_out0 = v_G2_12621_out0;
assign v_CARRY_5694_out0 = v_G2_13085_out0;
assign v_S_9231_out0 = v_G1_8085_out0;
assign v_S_9695_out0 = v_G1_8549_out0;
assign v_S_1396_out0 = v_S_9231_out0;
assign v_S_1620_out0 = v_S_9695_out0;
assign v_G1_4172_out0 = v_CARRY_5230_out0 || v_CARRY_5229_out0;
assign v_G1_4396_out0 = v_CARRY_5694_out0 || v_CARRY_5693_out0;
assign v_COUT_864_out0 = v_G1_4172_out0;
assign v_COUT_1088_out0 = v_G1_4396_out0;
assign v__4760_out0 = { v__7158_out0,v_S_1396_out0 };
assign v__4775_out0 = { v__7173_out0,v_S_1620_out0 };
assign v_CIN_9978_out0 = v_COUT_864_out0;
assign v_CIN_10202_out0 = v_COUT_1088_out0;
assign v_RD_6216_out0 = v_CIN_9978_out0;
assign v_RD_6680_out0 = v_CIN_10202_out0;
assign v_G1_8071_out0 = ((v_RD_6216_out0 && !v_RM_11656_out0) || (!v_RD_6216_out0) && v_RM_11656_out0);
assign v_G1_8535_out0 = ((v_RD_6680_out0 && !v_RM_12120_out0) || (!v_RD_6680_out0) && v_RM_12120_out0);
assign v_G2_12607_out0 = v_RD_6216_out0 && v_RM_11656_out0;
assign v_G2_13071_out0 = v_RD_6680_out0 && v_RM_12120_out0;
assign v_CARRY_5216_out0 = v_G2_12607_out0;
assign v_CARRY_5680_out0 = v_G2_13071_out0;
assign v_S_9217_out0 = v_G1_8071_out0;
assign v_S_9681_out0 = v_G1_8535_out0;
assign v_S_1389_out0 = v_S_9217_out0;
assign v_S_1613_out0 = v_S_9681_out0;
assign v_G1_4165_out0 = v_CARRY_5216_out0 || v_CARRY_5215_out0;
assign v_G1_4389_out0 = v_CARRY_5680_out0 || v_CARRY_5679_out0;
assign v_COUT_857_out0 = v_G1_4165_out0;
assign v_COUT_1081_out0 = v_G1_4389_out0;
assign v__6937_out0 = { v__4760_out0,v_S_1389_out0 };
assign v__6952_out0 = { v__4775_out0,v_S_1613_out0 };
assign v_CIN_9979_out0 = v_COUT_857_out0;
assign v_CIN_10203_out0 = v_COUT_1081_out0;
assign v_RD_6218_out0 = v_CIN_9979_out0;
assign v_RD_6682_out0 = v_CIN_10203_out0;
assign v_G1_8073_out0 = ((v_RD_6218_out0 && !v_RM_11658_out0) || (!v_RD_6218_out0) && v_RM_11658_out0);
assign v_G1_8537_out0 = ((v_RD_6682_out0 && !v_RM_12122_out0) || (!v_RD_6682_out0) && v_RM_12122_out0);
assign v_G2_12609_out0 = v_RD_6218_out0 && v_RM_11658_out0;
assign v_G2_13073_out0 = v_RD_6682_out0 && v_RM_12122_out0;
assign v_CARRY_5218_out0 = v_G2_12609_out0;
assign v_CARRY_5682_out0 = v_G2_13073_out0;
assign v_S_9219_out0 = v_G1_8073_out0;
assign v_S_9683_out0 = v_G1_8537_out0;
assign v_S_1390_out0 = v_S_9219_out0;
assign v_S_1614_out0 = v_S_9683_out0;
assign v_G1_4166_out0 = v_CARRY_5218_out0 || v_CARRY_5217_out0;
assign v_G1_4390_out0 = v_CARRY_5682_out0 || v_CARRY_5681_out0;
assign v_COUT_858_out0 = v_G1_4166_out0;
assign v_COUT_1082_out0 = v_G1_4390_out0;
assign v__5813_out0 = { v__6937_out0,v_S_1390_out0 };
assign v__5828_out0 = { v__6952_out0,v_S_1614_out0 };
assign v_CIN_9984_out0 = v_COUT_858_out0;
assign v_CIN_10208_out0 = v_COUT_1082_out0;
assign v_RD_6228_out0 = v_CIN_9984_out0;
assign v_RD_6692_out0 = v_CIN_10208_out0;
assign v_G1_8083_out0 = ((v_RD_6228_out0 && !v_RM_11668_out0) || (!v_RD_6228_out0) && v_RM_11668_out0);
assign v_G1_8547_out0 = ((v_RD_6692_out0 && !v_RM_12132_out0) || (!v_RD_6692_out0) && v_RM_12132_out0);
assign v_G2_12619_out0 = v_RD_6228_out0 && v_RM_11668_out0;
assign v_G2_13083_out0 = v_RD_6692_out0 && v_RM_12132_out0;
assign v_CARRY_5228_out0 = v_G2_12619_out0;
assign v_CARRY_5692_out0 = v_G2_13083_out0;
assign v_S_9229_out0 = v_G1_8083_out0;
assign v_S_9693_out0 = v_G1_8547_out0;
assign v_S_1395_out0 = v_S_9229_out0;
assign v_S_1619_out0 = v_S_9693_out0;
assign v_G1_4171_out0 = v_CARRY_5228_out0 || v_CARRY_5227_out0;
assign v_G1_4395_out0 = v_CARRY_5692_out0 || v_CARRY_5691_out0;
assign v_COUT_863_out0 = v_G1_4171_out0;
assign v_COUT_1087_out0 = v_G1_4395_out0;
assign v__2037_out0 = { v__5813_out0,v_S_1395_out0 };
assign v__2052_out0 = { v__5828_out0,v_S_1619_out0 };
assign v_CIN_9972_out0 = v_COUT_863_out0;
assign v_CIN_10196_out0 = v_COUT_1087_out0;
assign v_RD_6203_out0 = v_CIN_9972_out0;
assign v_RD_6667_out0 = v_CIN_10196_out0;
assign v_G1_8058_out0 = ((v_RD_6203_out0 && !v_RM_11643_out0) || (!v_RD_6203_out0) && v_RM_11643_out0);
assign v_G1_8522_out0 = ((v_RD_6667_out0 && !v_RM_12107_out0) || (!v_RD_6667_out0) && v_RM_12107_out0);
assign v_G2_12594_out0 = v_RD_6203_out0 && v_RM_11643_out0;
assign v_G2_13058_out0 = v_RD_6667_out0 && v_RM_12107_out0;
assign v_CARRY_5203_out0 = v_G2_12594_out0;
assign v_CARRY_5667_out0 = v_G2_13058_out0;
assign v_S_9204_out0 = v_G1_8058_out0;
assign v_S_9668_out0 = v_G1_8522_out0;
assign v_S_1383_out0 = v_S_9204_out0;
assign v_S_1607_out0 = v_S_9668_out0;
assign v_G1_4159_out0 = v_CARRY_5203_out0 || v_CARRY_5202_out0;
assign v_G1_4383_out0 = v_CARRY_5667_out0 || v_CARRY_5666_out0;
assign v_COUT_851_out0 = v_G1_4159_out0;
assign v_COUT_1075_out0 = v_G1_4383_out0;
assign v__2804_out0 = { v__2037_out0,v_S_1383_out0 };
assign v__2819_out0 = { v__2052_out0,v_S_1607_out0 };
assign v_CIN_9977_out0 = v_COUT_851_out0;
assign v_CIN_10201_out0 = v_COUT_1075_out0;
assign v_RD_6213_out0 = v_CIN_9977_out0;
assign v_RD_6677_out0 = v_CIN_10201_out0;
assign v_G1_8068_out0 = ((v_RD_6213_out0 && !v_RM_11653_out0) || (!v_RD_6213_out0) && v_RM_11653_out0);
assign v_G1_8532_out0 = ((v_RD_6677_out0 && !v_RM_12117_out0) || (!v_RD_6677_out0) && v_RM_12117_out0);
assign v_G2_12604_out0 = v_RD_6213_out0 && v_RM_11653_out0;
assign v_G2_13068_out0 = v_RD_6677_out0 && v_RM_12117_out0;
assign v_CARRY_5213_out0 = v_G2_12604_out0;
assign v_CARRY_5677_out0 = v_G2_13068_out0;
assign v_S_9214_out0 = v_G1_8068_out0;
assign v_S_9678_out0 = v_G1_8532_out0;
assign v_S_1388_out0 = v_S_9214_out0;
assign v_S_1612_out0 = v_S_9678_out0;
assign v_G1_4164_out0 = v_CARRY_5213_out0 || v_CARRY_5212_out0;
assign v_G1_4388_out0 = v_CARRY_5677_out0 || v_CARRY_5676_out0;
assign v_COUT_856_out0 = v_G1_4164_out0;
assign v_COUT_1080_out0 = v_G1_4388_out0;
assign v__1836_out0 = { v__2804_out0,v_S_1388_out0 };
assign v__1851_out0 = { v__2819_out0,v_S_1612_out0 };
assign v_CIN_9973_out0 = v_COUT_856_out0;
assign v_CIN_10197_out0 = v_COUT_1080_out0;
assign v_RD_6205_out0 = v_CIN_9973_out0;
assign v_RD_6669_out0 = v_CIN_10197_out0;
assign v_G1_8060_out0 = ((v_RD_6205_out0 && !v_RM_11645_out0) || (!v_RD_6205_out0) && v_RM_11645_out0);
assign v_G1_8524_out0 = ((v_RD_6669_out0 && !v_RM_12109_out0) || (!v_RD_6669_out0) && v_RM_12109_out0);
assign v_G2_12596_out0 = v_RD_6205_out0 && v_RM_11645_out0;
assign v_G2_13060_out0 = v_RD_6669_out0 && v_RM_12109_out0;
assign v_CARRY_5205_out0 = v_G2_12596_out0;
assign v_CARRY_5669_out0 = v_G2_13060_out0;
assign v_S_9206_out0 = v_G1_8060_out0;
assign v_S_9670_out0 = v_G1_8524_out0;
assign v_S_1384_out0 = v_S_9206_out0;
assign v_S_1608_out0 = v_S_9670_out0;
assign v_G1_4160_out0 = v_CARRY_5205_out0 || v_CARRY_5204_out0;
assign v_G1_4384_out0 = v_CARRY_5669_out0 || v_CARRY_5668_out0;
assign v_COUT_852_out0 = v_G1_4160_out0;
assign v_COUT_1076_out0 = v_G1_4384_out0;
assign v__4560_out0 = { v__1836_out0,v_S_1384_out0 };
assign v__4575_out0 = { v__1851_out0,v_S_1608_out0 };
assign v_RM_3521_out0 = v_COUT_852_out0;
assign v_RM_3745_out0 = v_COUT_1076_out0;
assign v_RM_11646_out0 = v_RM_3521_out0;
assign v_RM_12110_out0 = v_RM_3745_out0;
assign v_G1_8061_out0 = ((v_RD_6206_out0 && !v_RM_11646_out0) || (!v_RD_6206_out0) && v_RM_11646_out0);
assign v_G1_8525_out0 = ((v_RD_6670_out0 && !v_RM_12110_out0) || (!v_RD_6670_out0) && v_RM_12110_out0);
assign v_G2_12597_out0 = v_RD_6206_out0 && v_RM_11646_out0;
assign v_G2_13061_out0 = v_RD_6670_out0 && v_RM_12110_out0;
assign v_CARRY_5206_out0 = v_G2_12597_out0;
assign v_CARRY_5670_out0 = v_G2_13061_out0;
assign v_S_9207_out0 = v_G1_8061_out0;
assign v_S_9671_out0 = v_G1_8525_out0;
assign v_RM_11647_out0 = v_S_9207_out0;
assign v_RM_12111_out0 = v_S_9671_out0;
assign v_G1_8062_out0 = ((v_RD_6207_out0 && !v_RM_11647_out0) || (!v_RD_6207_out0) && v_RM_11647_out0);
assign v_G1_8526_out0 = ((v_RD_6671_out0 && !v_RM_12111_out0) || (!v_RD_6671_out0) && v_RM_12111_out0);
assign v_G2_12598_out0 = v_RD_6207_out0 && v_RM_11647_out0;
assign v_G2_13062_out0 = v_RD_6671_out0 && v_RM_12111_out0;
assign v_CARRY_5207_out0 = v_G2_12598_out0;
assign v_CARRY_5671_out0 = v_G2_13062_out0;
assign v_S_9208_out0 = v_G1_8062_out0;
assign v_S_9672_out0 = v_G1_8526_out0;
assign v_S_1385_out0 = v_S_9208_out0;
assign v_S_1609_out0 = v_S_9672_out0;
assign v_G1_4161_out0 = v_CARRY_5207_out0 || v_CARRY_5206_out0;
assign v_G1_4385_out0 = v_CARRY_5671_out0 || v_CARRY_5670_out0;
assign v_COUT_853_out0 = v_G1_4161_out0;
assign v_COUT_1077_out0 = v_G1_4385_out0;
assign v__10662_out0 = { v__4560_out0,v_S_1385_out0 };
assign v__10677_out0 = { v__4575_out0,v_S_1609_out0 };
assign v__10957_out0 = { v__10662_out0,v_COUT_853_out0 };
assign v__10972_out0 = { v__10677_out0,v_COUT_1077_out0 };
assign v_COUT_10927_out0 = v__10957_out0;
assign v_COUT_10942_out0 = v__10972_out0;
assign v_CIN_2364_out0 = v_COUT_10927_out0;
assign v_CIN_2379_out0 = v_COUT_10942_out0;
assign v__477_out0 = v_CIN_2364_out0[8:8];
assign v__492_out0 = v_CIN_2379_out0[8:8];
assign v__1782_out0 = v_CIN_2364_out0[6:6];
assign v__1797_out0 = v_CIN_2379_out0[6:6];
assign v__2164_out0 = v_CIN_2364_out0[3:3];
assign v__2179_out0 = v_CIN_2379_out0[3:3];
assign v__2203_out0 = v_CIN_2364_out0[15:15];
assign v__2217_out0 = v_CIN_2379_out0[15:15];
assign v__2511_out0 = v_CIN_2364_out0[0:0];
assign v__2526_out0 = v_CIN_2379_out0[0:0];
assign v__3060_out0 = v_CIN_2364_out0[9:9];
assign v__3075_out0 = v_CIN_2379_out0[9:9];
assign v__3094_out0 = v_CIN_2364_out0[2:2];
assign v__3109_out0 = v_CIN_2379_out0[2:2];
assign v__3148_out0 = v_CIN_2364_out0[7:7];
assign v__3163_out0 = v_CIN_2379_out0[7:7];
assign v__3832_out0 = v_CIN_2364_out0[1:1];
assign v__3847_out0 = v_CIN_2379_out0[1:1];
assign v__3870_out0 = v_CIN_2364_out0[10:10];
assign v__3885_out0 = v_CIN_2379_out0[10:10];
assign v__6809_out0 = v_CIN_2364_out0[11:11];
assign v__6824_out0 = v_CIN_2379_out0[11:11];
assign v__7653_out0 = v_CIN_2364_out0[12:12];
assign v__7668_out0 = v_CIN_2379_out0[12:12];
assign v__8708_out0 = v_CIN_2364_out0[13:13];
assign v__8723_out0 = v_CIN_2379_out0[13:13];
assign v__8778_out0 = v_CIN_2364_out0[14:14];
assign v__8793_out0 = v_CIN_2379_out0[14:14];
assign v__10728_out0 = v_CIN_2364_out0[5:5];
assign v__10743_out0 = v_CIN_2379_out0[5:5];
assign v__13457_out0 = v_CIN_2364_out0[4:4];
assign v__13472_out0 = v_CIN_2379_out0[4:4];
assign v_RM_3489_out0 = v__7653_out0;
assign v_RM_3490_out0 = v__8778_out0;
assign v_RM_3492_out0 = v__10728_out0;
assign v_RM_3493_out0 = v__13457_out0;
assign v_RM_3494_out0 = v__8708_out0;
assign v_RM_3495_out0 = v__3060_out0;
assign v_RM_3496_out0 = v__3870_out0;
assign v_RM_3497_out0 = v__3832_out0;
assign v_RM_3498_out0 = v__2164_out0;
assign v_RM_3499_out0 = v__1782_out0;
assign v_RM_3500_out0 = v__3148_out0;
assign v_RM_3501_out0 = v__6809_out0;
assign v_RM_3502_out0 = v__477_out0;
assign v_RM_3503_out0 = v__3094_out0;
assign v_RM_3713_out0 = v__7668_out0;
assign v_RM_3714_out0 = v__8793_out0;
assign v_RM_3716_out0 = v__10743_out0;
assign v_RM_3717_out0 = v__13472_out0;
assign v_RM_3718_out0 = v__8723_out0;
assign v_RM_3719_out0 = v__3075_out0;
assign v_RM_3720_out0 = v__3885_out0;
assign v_RM_3721_out0 = v__3847_out0;
assign v_RM_3722_out0 = v__2179_out0;
assign v_RM_3723_out0 = v__1797_out0;
assign v_RM_3724_out0 = v__3163_out0;
assign v_RM_3725_out0 = v__6824_out0;
assign v_RM_3726_out0 = v__492_out0;
assign v_RM_3727_out0 = v__3109_out0;
assign v_CIN_9944_out0 = v__2203_out0;
assign v_CIN_10168_out0 = v__2217_out0;
assign v_RM_11592_out0 = v__2511_out0;
assign v_RM_12056_out0 = v__2526_out0;
assign v_RD_6145_out0 = v_CIN_9944_out0;
assign v_RD_6609_out0 = v_CIN_10168_out0;
assign v_G1_8007_out0 = ((v_RD_6152_out0 && !v_RM_11592_out0) || (!v_RD_6152_out0) && v_RM_11592_out0);
assign v_G1_8471_out0 = ((v_RD_6616_out0 && !v_RM_12056_out0) || (!v_RD_6616_out0) && v_RM_12056_out0);
assign v_RM_11580_out0 = v_RM_3489_out0;
assign v_RM_11582_out0 = v_RM_3490_out0;
assign v_RM_11586_out0 = v_RM_3492_out0;
assign v_RM_11588_out0 = v_RM_3493_out0;
assign v_RM_11590_out0 = v_RM_3494_out0;
assign v_RM_11593_out0 = v_RM_3495_out0;
assign v_RM_11595_out0 = v_RM_3496_out0;
assign v_RM_11597_out0 = v_RM_3497_out0;
assign v_RM_11599_out0 = v_RM_3498_out0;
assign v_RM_11601_out0 = v_RM_3499_out0;
assign v_RM_11603_out0 = v_RM_3500_out0;
assign v_RM_11605_out0 = v_RM_3501_out0;
assign v_RM_11607_out0 = v_RM_3502_out0;
assign v_RM_11609_out0 = v_RM_3503_out0;
assign v_RM_12044_out0 = v_RM_3713_out0;
assign v_RM_12046_out0 = v_RM_3714_out0;
assign v_RM_12050_out0 = v_RM_3716_out0;
assign v_RM_12052_out0 = v_RM_3717_out0;
assign v_RM_12054_out0 = v_RM_3718_out0;
assign v_RM_12057_out0 = v_RM_3719_out0;
assign v_RM_12059_out0 = v_RM_3720_out0;
assign v_RM_12061_out0 = v_RM_3721_out0;
assign v_RM_12063_out0 = v_RM_3722_out0;
assign v_RM_12065_out0 = v_RM_3723_out0;
assign v_RM_12067_out0 = v_RM_3724_out0;
assign v_RM_12069_out0 = v_RM_3725_out0;
assign v_RM_12071_out0 = v_RM_3726_out0;
assign v_RM_12073_out0 = v_RM_3727_out0;
assign v_G2_12543_out0 = v_RD_6152_out0 && v_RM_11592_out0;
assign v_G2_13007_out0 = v_RD_6616_out0 && v_RM_12056_out0;
assign v_CARRY_5152_out0 = v_G2_12543_out0;
assign v_CARRY_5616_out0 = v_G2_13007_out0;
assign v_G1_7995_out0 = ((v_RD_6140_out0 && !v_RM_11580_out0) || (!v_RD_6140_out0) && v_RM_11580_out0);
assign v_G1_7997_out0 = ((v_RD_6142_out0 && !v_RM_11582_out0) || (!v_RD_6142_out0) && v_RM_11582_out0);
assign v_G1_8001_out0 = ((v_RD_6146_out0 && !v_RM_11586_out0) || (!v_RD_6146_out0) && v_RM_11586_out0);
assign v_G1_8003_out0 = ((v_RD_6148_out0 && !v_RM_11588_out0) || (!v_RD_6148_out0) && v_RM_11588_out0);
assign v_G1_8005_out0 = ((v_RD_6150_out0 && !v_RM_11590_out0) || (!v_RD_6150_out0) && v_RM_11590_out0);
assign v_G1_8008_out0 = ((v_RD_6153_out0 && !v_RM_11593_out0) || (!v_RD_6153_out0) && v_RM_11593_out0);
assign v_G1_8010_out0 = ((v_RD_6155_out0 && !v_RM_11595_out0) || (!v_RD_6155_out0) && v_RM_11595_out0);
assign v_G1_8012_out0 = ((v_RD_6157_out0 && !v_RM_11597_out0) || (!v_RD_6157_out0) && v_RM_11597_out0);
assign v_G1_8014_out0 = ((v_RD_6159_out0 && !v_RM_11599_out0) || (!v_RD_6159_out0) && v_RM_11599_out0);
assign v_G1_8016_out0 = ((v_RD_6161_out0 && !v_RM_11601_out0) || (!v_RD_6161_out0) && v_RM_11601_out0);
assign v_G1_8018_out0 = ((v_RD_6163_out0 && !v_RM_11603_out0) || (!v_RD_6163_out0) && v_RM_11603_out0);
assign v_G1_8020_out0 = ((v_RD_6165_out0 && !v_RM_11605_out0) || (!v_RD_6165_out0) && v_RM_11605_out0);
assign v_G1_8022_out0 = ((v_RD_6167_out0 && !v_RM_11607_out0) || (!v_RD_6167_out0) && v_RM_11607_out0);
assign v_G1_8024_out0 = ((v_RD_6169_out0 && !v_RM_11609_out0) || (!v_RD_6169_out0) && v_RM_11609_out0);
assign v_G1_8459_out0 = ((v_RD_6604_out0 && !v_RM_12044_out0) || (!v_RD_6604_out0) && v_RM_12044_out0);
assign v_G1_8461_out0 = ((v_RD_6606_out0 && !v_RM_12046_out0) || (!v_RD_6606_out0) && v_RM_12046_out0);
assign v_G1_8465_out0 = ((v_RD_6610_out0 && !v_RM_12050_out0) || (!v_RD_6610_out0) && v_RM_12050_out0);
assign v_G1_8467_out0 = ((v_RD_6612_out0 && !v_RM_12052_out0) || (!v_RD_6612_out0) && v_RM_12052_out0);
assign v_G1_8469_out0 = ((v_RD_6614_out0 && !v_RM_12054_out0) || (!v_RD_6614_out0) && v_RM_12054_out0);
assign v_G1_8472_out0 = ((v_RD_6617_out0 && !v_RM_12057_out0) || (!v_RD_6617_out0) && v_RM_12057_out0);
assign v_G1_8474_out0 = ((v_RD_6619_out0 && !v_RM_12059_out0) || (!v_RD_6619_out0) && v_RM_12059_out0);
assign v_G1_8476_out0 = ((v_RD_6621_out0 && !v_RM_12061_out0) || (!v_RD_6621_out0) && v_RM_12061_out0);
assign v_G1_8478_out0 = ((v_RD_6623_out0 && !v_RM_12063_out0) || (!v_RD_6623_out0) && v_RM_12063_out0);
assign v_G1_8480_out0 = ((v_RD_6625_out0 && !v_RM_12065_out0) || (!v_RD_6625_out0) && v_RM_12065_out0);
assign v_G1_8482_out0 = ((v_RD_6627_out0 && !v_RM_12067_out0) || (!v_RD_6627_out0) && v_RM_12067_out0);
assign v_G1_8484_out0 = ((v_RD_6629_out0 && !v_RM_12069_out0) || (!v_RD_6629_out0) && v_RM_12069_out0);
assign v_G1_8486_out0 = ((v_RD_6631_out0 && !v_RM_12071_out0) || (!v_RD_6631_out0) && v_RM_12071_out0);
assign v_G1_8488_out0 = ((v_RD_6633_out0 && !v_RM_12073_out0) || (!v_RD_6633_out0) && v_RM_12073_out0);
assign v_S_9153_out0 = v_G1_8007_out0;
assign v_S_9617_out0 = v_G1_8471_out0;
assign v_G2_12531_out0 = v_RD_6140_out0 && v_RM_11580_out0;
assign v_G2_12533_out0 = v_RD_6142_out0 && v_RM_11582_out0;
assign v_G2_12537_out0 = v_RD_6146_out0 && v_RM_11586_out0;
assign v_G2_12539_out0 = v_RD_6148_out0 && v_RM_11588_out0;
assign v_G2_12541_out0 = v_RD_6150_out0 && v_RM_11590_out0;
assign v_G2_12544_out0 = v_RD_6153_out0 && v_RM_11593_out0;
assign v_G2_12546_out0 = v_RD_6155_out0 && v_RM_11595_out0;
assign v_G2_12548_out0 = v_RD_6157_out0 && v_RM_11597_out0;
assign v_G2_12550_out0 = v_RD_6159_out0 && v_RM_11599_out0;
assign v_G2_12552_out0 = v_RD_6161_out0 && v_RM_11601_out0;
assign v_G2_12554_out0 = v_RD_6163_out0 && v_RM_11603_out0;
assign v_G2_12556_out0 = v_RD_6165_out0 && v_RM_11605_out0;
assign v_G2_12558_out0 = v_RD_6167_out0 && v_RM_11607_out0;
assign v_G2_12560_out0 = v_RD_6169_out0 && v_RM_11609_out0;
assign v_G2_12995_out0 = v_RD_6604_out0 && v_RM_12044_out0;
assign v_G2_12997_out0 = v_RD_6606_out0 && v_RM_12046_out0;
assign v_G2_13001_out0 = v_RD_6610_out0 && v_RM_12050_out0;
assign v_G2_13003_out0 = v_RD_6612_out0 && v_RM_12052_out0;
assign v_G2_13005_out0 = v_RD_6614_out0 && v_RM_12054_out0;
assign v_G2_13008_out0 = v_RD_6617_out0 && v_RM_12057_out0;
assign v_G2_13010_out0 = v_RD_6619_out0 && v_RM_12059_out0;
assign v_G2_13012_out0 = v_RD_6621_out0 && v_RM_12061_out0;
assign v_G2_13014_out0 = v_RD_6623_out0 && v_RM_12063_out0;
assign v_G2_13016_out0 = v_RD_6625_out0 && v_RM_12065_out0;
assign v_G2_13018_out0 = v_RD_6627_out0 && v_RM_12067_out0;
assign v_G2_13020_out0 = v_RD_6629_out0 && v_RM_12069_out0;
assign v_G2_13022_out0 = v_RD_6631_out0 && v_RM_12071_out0;
assign v_G2_13024_out0 = v_RD_6633_out0 && v_RM_12073_out0;
assign v_S_4674_out0 = v_S_9153_out0;
assign v_S_4689_out0 = v_S_9617_out0;
assign v_CARRY_5140_out0 = v_G2_12531_out0;
assign v_CARRY_5142_out0 = v_G2_12533_out0;
assign v_CARRY_5146_out0 = v_G2_12537_out0;
assign v_CARRY_5148_out0 = v_G2_12539_out0;
assign v_CARRY_5150_out0 = v_G2_12541_out0;
assign v_CARRY_5153_out0 = v_G2_12544_out0;
assign v_CARRY_5155_out0 = v_G2_12546_out0;
assign v_CARRY_5157_out0 = v_G2_12548_out0;
assign v_CARRY_5159_out0 = v_G2_12550_out0;
assign v_CARRY_5161_out0 = v_G2_12552_out0;
assign v_CARRY_5163_out0 = v_G2_12554_out0;
assign v_CARRY_5165_out0 = v_G2_12556_out0;
assign v_CARRY_5167_out0 = v_G2_12558_out0;
assign v_CARRY_5169_out0 = v_G2_12560_out0;
assign v_CARRY_5604_out0 = v_G2_12995_out0;
assign v_CARRY_5606_out0 = v_G2_12997_out0;
assign v_CARRY_5610_out0 = v_G2_13001_out0;
assign v_CARRY_5612_out0 = v_G2_13003_out0;
assign v_CARRY_5614_out0 = v_G2_13005_out0;
assign v_CARRY_5617_out0 = v_G2_13008_out0;
assign v_CARRY_5619_out0 = v_G2_13010_out0;
assign v_CARRY_5621_out0 = v_G2_13012_out0;
assign v_CARRY_5623_out0 = v_G2_13014_out0;
assign v_CARRY_5625_out0 = v_G2_13016_out0;
assign v_CARRY_5627_out0 = v_G2_13018_out0;
assign v_CARRY_5629_out0 = v_G2_13020_out0;
assign v_CARRY_5631_out0 = v_G2_13022_out0;
assign v_CARRY_5633_out0 = v_G2_13024_out0;
assign v_S_9141_out0 = v_G1_7995_out0;
assign v_S_9143_out0 = v_G1_7997_out0;
assign v_S_9147_out0 = v_G1_8001_out0;
assign v_S_9149_out0 = v_G1_8003_out0;
assign v_S_9151_out0 = v_G1_8005_out0;
assign v_S_9154_out0 = v_G1_8008_out0;
assign v_S_9156_out0 = v_G1_8010_out0;
assign v_S_9158_out0 = v_G1_8012_out0;
assign v_S_9160_out0 = v_G1_8014_out0;
assign v_S_9162_out0 = v_G1_8016_out0;
assign v_S_9164_out0 = v_G1_8018_out0;
assign v_S_9166_out0 = v_G1_8020_out0;
assign v_S_9168_out0 = v_G1_8022_out0;
assign v_S_9170_out0 = v_G1_8024_out0;
assign v_S_9605_out0 = v_G1_8459_out0;
assign v_S_9607_out0 = v_G1_8461_out0;
assign v_S_9611_out0 = v_G1_8465_out0;
assign v_S_9613_out0 = v_G1_8467_out0;
assign v_S_9615_out0 = v_G1_8469_out0;
assign v_S_9618_out0 = v_G1_8472_out0;
assign v_S_9620_out0 = v_G1_8474_out0;
assign v_S_9622_out0 = v_G1_8476_out0;
assign v_S_9624_out0 = v_G1_8478_out0;
assign v_S_9626_out0 = v_G1_8480_out0;
assign v_S_9628_out0 = v_G1_8482_out0;
assign v_S_9630_out0 = v_G1_8484_out0;
assign v_S_9632_out0 = v_G1_8486_out0;
assign v_S_9634_out0 = v_G1_8488_out0;
assign v_CIN_9950_out0 = v_CARRY_5152_out0;
assign v_CIN_10174_out0 = v_CARRY_5616_out0;
assign v__43_out0 = { v__636_out0,v_S_4674_out0 };
assign v__44_out0 = { v__637_out0,v_S_4689_out0 };
assign v_RD_6158_out0 = v_CIN_9950_out0;
assign v_RD_6622_out0 = v_CIN_10174_out0;
assign v_RM_11581_out0 = v_S_9141_out0;
assign v_RM_11583_out0 = v_S_9143_out0;
assign v_RM_11587_out0 = v_S_9147_out0;
assign v_RM_11589_out0 = v_S_9149_out0;
assign v_RM_11591_out0 = v_S_9151_out0;
assign v_RM_11594_out0 = v_S_9154_out0;
assign v_RM_11596_out0 = v_S_9156_out0;
assign v_RM_11598_out0 = v_S_9158_out0;
assign v_RM_11600_out0 = v_S_9160_out0;
assign v_RM_11602_out0 = v_S_9162_out0;
assign v_RM_11604_out0 = v_S_9164_out0;
assign v_RM_11606_out0 = v_S_9166_out0;
assign v_RM_11608_out0 = v_S_9168_out0;
assign v_RM_11610_out0 = v_S_9170_out0;
assign v_RM_12045_out0 = v_S_9605_out0;
assign v_RM_12047_out0 = v_S_9607_out0;
assign v_RM_12051_out0 = v_S_9611_out0;
assign v_RM_12053_out0 = v_S_9613_out0;
assign v_RM_12055_out0 = v_S_9615_out0;
assign v_RM_12058_out0 = v_S_9618_out0;
assign v_RM_12060_out0 = v_S_9620_out0;
assign v_RM_12062_out0 = v_S_9622_out0;
assign v_RM_12064_out0 = v_S_9624_out0;
assign v_RM_12066_out0 = v_S_9626_out0;
assign v_RM_12068_out0 = v_S_9628_out0;
assign v_RM_12070_out0 = v_S_9630_out0;
assign v_RM_12072_out0 = v_S_9632_out0;
assign v_RM_12074_out0 = v_S_9634_out0;
assign v_G1_8013_out0 = ((v_RD_6158_out0 && !v_RM_11598_out0) || (!v_RD_6158_out0) && v_RM_11598_out0);
assign v_G1_8477_out0 = ((v_RD_6622_out0 && !v_RM_12062_out0) || (!v_RD_6622_out0) && v_RM_12062_out0);
assign v_G2_12549_out0 = v_RD_6158_out0 && v_RM_11598_out0;
assign v_G2_13013_out0 = v_RD_6622_out0 && v_RM_12062_out0;
assign v_CARRY_5158_out0 = v_G2_12549_out0;
assign v_CARRY_5622_out0 = v_G2_13013_out0;
assign v_S_9159_out0 = v_G1_8013_out0;
assign v_S_9623_out0 = v_G1_8477_out0;
assign v_S_1361_out0 = v_S_9159_out0;
assign v_S_1585_out0 = v_S_9623_out0;
assign v_G1_4137_out0 = v_CARRY_5158_out0 || v_CARRY_5157_out0;
assign v_G1_4361_out0 = v_CARRY_5622_out0 || v_CARRY_5621_out0;
assign v_COUT_829_out0 = v_G1_4137_out0;
assign v_COUT_1053_out0 = v_G1_4361_out0;
assign v_CIN_9956_out0 = v_COUT_829_out0;
assign v_CIN_10180_out0 = v_COUT_1053_out0;
assign v_RD_6170_out0 = v_CIN_9956_out0;
assign v_RD_6634_out0 = v_CIN_10180_out0;
assign v_G1_8025_out0 = ((v_RD_6170_out0 && !v_RM_11610_out0) || (!v_RD_6170_out0) && v_RM_11610_out0);
assign v_G1_8489_out0 = ((v_RD_6634_out0 && !v_RM_12074_out0) || (!v_RD_6634_out0) && v_RM_12074_out0);
assign v_G2_12561_out0 = v_RD_6170_out0 && v_RM_11610_out0;
assign v_G2_13025_out0 = v_RD_6634_out0 && v_RM_12074_out0;
assign v_CARRY_5170_out0 = v_G2_12561_out0;
assign v_CARRY_5634_out0 = v_G2_13025_out0;
assign v_S_9171_out0 = v_G1_8025_out0;
assign v_S_9635_out0 = v_G1_8489_out0;
assign v_S_1367_out0 = v_S_9171_out0;
assign v_S_1591_out0 = v_S_9635_out0;
assign v_G1_4143_out0 = v_CARRY_5170_out0 || v_CARRY_5169_out0;
assign v_G1_4367_out0 = v_CARRY_5634_out0 || v_CARRY_5633_out0;
assign v_COUT_835_out0 = v_G1_4143_out0;
assign v_COUT_1059_out0 = v_G1_4367_out0;
assign v__4791_out0 = { v_S_1361_out0,v_S_1367_out0 };
assign v__4806_out0 = { v_S_1585_out0,v_S_1591_out0 };
assign v_CIN_9951_out0 = v_COUT_835_out0;
assign v_CIN_10175_out0 = v_COUT_1059_out0;
assign v_RD_6160_out0 = v_CIN_9951_out0;
assign v_RD_6624_out0 = v_CIN_10175_out0;
assign v_G1_8015_out0 = ((v_RD_6160_out0 && !v_RM_11600_out0) || (!v_RD_6160_out0) && v_RM_11600_out0);
assign v_G1_8479_out0 = ((v_RD_6624_out0 && !v_RM_12064_out0) || (!v_RD_6624_out0) && v_RM_12064_out0);
assign v_G2_12551_out0 = v_RD_6160_out0 && v_RM_11600_out0;
assign v_G2_13015_out0 = v_RD_6624_out0 && v_RM_12064_out0;
assign v_CARRY_5160_out0 = v_G2_12551_out0;
assign v_CARRY_5624_out0 = v_G2_13015_out0;
assign v_S_9161_out0 = v_G1_8015_out0;
assign v_S_9625_out0 = v_G1_8479_out0;
assign v_S_1362_out0 = v_S_9161_out0;
assign v_S_1586_out0 = v_S_9625_out0;
assign v_G1_4138_out0 = v_CARRY_5160_out0 || v_CARRY_5159_out0;
assign v_G1_4362_out0 = v_CARRY_5624_out0 || v_CARRY_5623_out0;
assign v_COUT_830_out0 = v_G1_4138_out0;
assign v_COUT_1054_out0 = v_G1_4362_out0;
assign v__2561_out0 = { v__4791_out0,v_S_1362_out0 };
assign v__2576_out0 = { v__4806_out0,v_S_1586_out0 };
assign v_CIN_9946_out0 = v_COUT_830_out0;
assign v_CIN_10170_out0 = v_COUT_1054_out0;
assign v_RD_6149_out0 = v_CIN_9946_out0;
assign v_RD_6613_out0 = v_CIN_10170_out0;
assign v_G1_8004_out0 = ((v_RD_6149_out0 && !v_RM_11589_out0) || (!v_RD_6149_out0) && v_RM_11589_out0);
assign v_G1_8468_out0 = ((v_RD_6613_out0 && !v_RM_12053_out0) || (!v_RD_6613_out0) && v_RM_12053_out0);
assign v_G2_12540_out0 = v_RD_6149_out0 && v_RM_11589_out0;
assign v_G2_13004_out0 = v_RD_6613_out0 && v_RM_12053_out0;
assign v_CARRY_5149_out0 = v_G2_12540_out0;
assign v_CARRY_5613_out0 = v_G2_13004_out0;
assign v_S_9150_out0 = v_G1_8004_out0;
assign v_S_9614_out0 = v_G1_8468_out0;
assign v_S_1357_out0 = v_S_9150_out0;
assign v_S_1581_out0 = v_S_9614_out0;
assign v_G1_4133_out0 = v_CARRY_5149_out0 || v_CARRY_5148_out0;
assign v_G1_4357_out0 = v_CARRY_5613_out0 || v_CARRY_5612_out0;
assign v_COUT_825_out0 = v_G1_4133_out0;
assign v_COUT_1049_out0 = v_G1_4357_out0;
assign v__7041_out0 = { v__2561_out0,v_S_1357_out0 };
assign v__7056_out0 = { v__2576_out0,v_S_1581_out0 };
assign v_CIN_9945_out0 = v_COUT_825_out0;
assign v_CIN_10169_out0 = v_COUT_1049_out0;
assign v_RD_6147_out0 = v_CIN_9945_out0;
assign v_RD_6611_out0 = v_CIN_10169_out0;
assign v_G1_8002_out0 = ((v_RD_6147_out0 && !v_RM_11587_out0) || (!v_RD_6147_out0) && v_RM_11587_out0);
assign v_G1_8466_out0 = ((v_RD_6611_out0 && !v_RM_12051_out0) || (!v_RD_6611_out0) && v_RM_12051_out0);
assign v_G2_12538_out0 = v_RD_6147_out0 && v_RM_11587_out0;
assign v_G2_13002_out0 = v_RD_6611_out0 && v_RM_12051_out0;
assign v_CARRY_5147_out0 = v_G2_12538_out0;
assign v_CARRY_5611_out0 = v_G2_13002_out0;
assign v_S_9148_out0 = v_G1_8002_out0;
assign v_S_9612_out0 = v_G1_8466_out0;
assign v_S_1356_out0 = v_S_9148_out0;
assign v_S_1580_out0 = v_S_9612_out0;
assign v_G1_4132_out0 = v_CARRY_5147_out0 || v_CARRY_5146_out0;
assign v_G1_4356_out0 = v_CARRY_5611_out0 || v_CARRY_5610_out0;
assign v_COUT_824_out0 = v_G1_4132_out0;
assign v_COUT_1048_out0 = v_G1_4356_out0;
assign v__13527_out0 = { v__7041_out0,v_S_1356_out0 };
assign v__13542_out0 = { v__7056_out0,v_S_1580_out0 };
assign v_CIN_9952_out0 = v_COUT_824_out0;
assign v_CIN_10176_out0 = v_COUT_1048_out0;
assign v_RD_6162_out0 = v_CIN_9952_out0;
assign v_RD_6626_out0 = v_CIN_10176_out0;
assign v_G1_8017_out0 = ((v_RD_6162_out0 && !v_RM_11602_out0) || (!v_RD_6162_out0) && v_RM_11602_out0);
assign v_G1_8481_out0 = ((v_RD_6626_out0 && !v_RM_12066_out0) || (!v_RD_6626_out0) && v_RM_12066_out0);
assign v_G2_12553_out0 = v_RD_6162_out0 && v_RM_11602_out0;
assign v_G2_13017_out0 = v_RD_6626_out0 && v_RM_12066_out0;
assign v_CARRY_5162_out0 = v_G2_12553_out0;
assign v_CARRY_5626_out0 = v_G2_13017_out0;
assign v_S_9163_out0 = v_G1_8017_out0;
assign v_S_9627_out0 = v_G1_8481_out0;
assign v_S_1363_out0 = v_S_9163_out0;
assign v_S_1587_out0 = v_S_9627_out0;
assign v_G1_4139_out0 = v_CARRY_5162_out0 || v_CARRY_5161_out0;
assign v_G1_4363_out0 = v_CARRY_5626_out0 || v_CARRY_5625_out0;
assign v_COUT_831_out0 = v_G1_4139_out0;
assign v_COUT_1055_out0 = v_G1_4363_out0;
assign v__3320_out0 = { v__13527_out0,v_S_1363_out0 };
assign v__3335_out0 = { v__13542_out0,v_S_1587_out0 };
assign v_CIN_9953_out0 = v_COUT_831_out0;
assign v_CIN_10177_out0 = v_COUT_1055_out0;
assign v_RD_6164_out0 = v_CIN_9953_out0;
assign v_RD_6628_out0 = v_CIN_10177_out0;
assign v_G1_8019_out0 = ((v_RD_6164_out0 && !v_RM_11604_out0) || (!v_RD_6164_out0) && v_RM_11604_out0);
assign v_G1_8483_out0 = ((v_RD_6628_out0 && !v_RM_12068_out0) || (!v_RD_6628_out0) && v_RM_12068_out0);
assign v_G2_12555_out0 = v_RD_6164_out0 && v_RM_11604_out0;
assign v_G2_13019_out0 = v_RD_6628_out0 && v_RM_12068_out0;
assign v_CARRY_5164_out0 = v_G2_12555_out0;
assign v_CARRY_5628_out0 = v_G2_13019_out0;
assign v_S_9165_out0 = v_G1_8019_out0;
assign v_S_9629_out0 = v_G1_8483_out0;
assign v_S_1364_out0 = v_S_9165_out0;
assign v_S_1588_out0 = v_S_9629_out0;
assign v_G1_4140_out0 = v_CARRY_5164_out0 || v_CARRY_5163_out0;
assign v_G1_4364_out0 = v_CARRY_5628_out0 || v_CARRY_5627_out0;
assign v_COUT_832_out0 = v_G1_4140_out0;
assign v_COUT_1056_out0 = v_G1_4364_out0;
assign v__7156_out0 = { v__3320_out0,v_S_1364_out0 };
assign v__7171_out0 = { v__3335_out0,v_S_1588_out0 };
assign v_CIN_9955_out0 = v_COUT_832_out0;
assign v_CIN_10179_out0 = v_COUT_1056_out0;
assign v_RD_6168_out0 = v_CIN_9955_out0;
assign v_RD_6632_out0 = v_CIN_10179_out0;
assign v_G1_8023_out0 = ((v_RD_6168_out0 && !v_RM_11608_out0) || (!v_RD_6168_out0) && v_RM_11608_out0);
assign v_G1_8487_out0 = ((v_RD_6632_out0 && !v_RM_12072_out0) || (!v_RD_6632_out0) && v_RM_12072_out0);
assign v_G2_12559_out0 = v_RD_6168_out0 && v_RM_11608_out0;
assign v_G2_13023_out0 = v_RD_6632_out0 && v_RM_12072_out0;
assign v_CARRY_5168_out0 = v_G2_12559_out0;
assign v_CARRY_5632_out0 = v_G2_13023_out0;
assign v_S_9169_out0 = v_G1_8023_out0;
assign v_S_9633_out0 = v_G1_8487_out0;
assign v_S_1366_out0 = v_S_9169_out0;
assign v_S_1590_out0 = v_S_9633_out0;
assign v_G1_4142_out0 = v_CARRY_5168_out0 || v_CARRY_5167_out0;
assign v_G1_4366_out0 = v_CARRY_5632_out0 || v_CARRY_5631_out0;
assign v_COUT_834_out0 = v_G1_4142_out0;
assign v_COUT_1058_out0 = v_G1_4366_out0;
assign v__4758_out0 = { v__7156_out0,v_S_1366_out0 };
assign v__4773_out0 = { v__7171_out0,v_S_1590_out0 };
assign v_CIN_9948_out0 = v_COUT_834_out0;
assign v_CIN_10172_out0 = v_COUT_1058_out0;
assign v_RD_6154_out0 = v_CIN_9948_out0;
assign v_RD_6618_out0 = v_CIN_10172_out0;
assign v_G1_8009_out0 = ((v_RD_6154_out0 && !v_RM_11594_out0) || (!v_RD_6154_out0) && v_RM_11594_out0);
assign v_G1_8473_out0 = ((v_RD_6618_out0 && !v_RM_12058_out0) || (!v_RD_6618_out0) && v_RM_12058_out0);
assign v_G2_12545_out0 = v_RD_6154_out0 && v_RM_11594_out0;
assign v_G2_13009_out0 = v_RD_6618_out0 && v_RM_12058_out0;
assign v_CARRY_5154_out0 = v_G2_12545_out0;
assign v_CARRY_5618_out0 = v_G2_13009_out0;
assign v_S_9155_out0 = v_G1_8009_out0;
assign v_S_9619_out0 = v_G1_8473_out0;
assign v_S_1359_out0 = v_S_9155_out0;
assign v_S_1583_out0 = v_S_9619_out0;
assign v_G1_4135_out0 = v_CARRY_5154_out0 || v_CARRY_5153_out0;
assign v_G1_4359_out0 = v_CARRY_5618_out0 || v_CARRY_5617_out0;
assign v_COUT_827_out0 = v_G1_4135_out0;
assign v_COUT_1051_out0 = v_G1_4359_out0;
assign v__6935_out0 = { v__4758_out0,v_S_1359_out0 };
assign v__6950_out0 = { v__4773_out0,v_S_1583_out0 };
assign v_CIN_9949_out0 = v_COUT_827_out0;
assign v_CIN_10173_out0 = v_COUT_1051_out0;
assign v_RD_6156_out0 = v_CIN_9949_out0;
assign v_RD_6620_out0 = v_CIN_10173_out0;
assign v_G1_8011_out0 = ((v_RD_6156_out0 && !v_RM_11596_out0) || (!v_RD_6156_out0) && v_RM_11596_out0);
assign v_G1_8475_out0 = ((v_RD_6620_out0 && !v_RM_12060_out0) || (!v_RD_6620_out0) && v_RM_12060_out0);
assign v_G2_12547_out0 = v_RD_6156_out0 && v_RM_11596_out0;
assign v_G2_13011_out0 = v_RD_6620_out0 && v_RM_12060_out0;
assign v_CARRY_5156_out0 = v_G2_12547_out0;
assign v_CARRY_5620_out0 = v_G2_13011_out0;
assign v_S_9157_out0 = v_G1_8011_out0;
assign v_S_9621_out0 = v_G1_8475_out0;
assign v_S_1360_out0 = v_S_9157_out0;
assign v_S_1584_out0 = v_S_9621_out0;
assign v_G1_4136_out0 = v_CARRY_5156_out0 || v_CARRY_5155_out0;
assign v_G1_4360_out0 = v_CARRY_5620_out0 || v_CARRY_5619_out0;
assign v_COUT_828_out0 = v_G1_4136_out0;
assign v_COUT_1052_out0 = v_G1_4360_out0;
assign v__5811_out0 = { v__6935_out0,v_S_1360_out0 };
assign v__5826_out0 = { v__6950_out0,v_S_1584_out0 };
assign v_CIN_9954_out0 = v_COUT_828_out0;
assign v_CIN_10178_out0 = v_COUT_1052_out0;
assign v_RD_6166_out0 = v_CIN_9954_out0;
assign v_RD_6630_out0 = v_CIN_10178_out0;
assign v_G1_8021_out0 = ((v_RD_6166_out0 && !v_RM_11606_out0) || (!v_RD_6166_out0) && v_RM_11606_out0);
assign v_G1_8485_out0 = ((v_RD_6630_out0 && !v_RM_12070_out0) || (!v_RD_6630_out0) && v_RM_12070_out0);
assign v_G2_12557_out0 = v_RD_6166_out0 && v_RM_11606_out0;
assign v_G2_13021_out0 = v_RD_6630_out0 && v_RM_12070_out0;
assign v_CARRY_5166_out0 = v_G2_12557_out0;
assign v_CARRY_5630_out0 = v_G2_13021_out0;
assign v_S_9167_out0 = v_G1_8021_out0;
assign v_S_9631_out0 = v_G1_8485_out0;
assign v_S_1365_out0 = v_S_9167_out0;
assign v_S_1589_out0 = v_S_9631_out0;
assign v_G1_4141_out0 = v_CARRY_5166_out0 || v_CARRY_5165_out0;
assign v_G1_4365_out0 = v_CARRY_5630_out0 || v_CARRY_5629_out0;
assign v_COUT_833_out0 = v_G1_4141_out0;
assign v_COUT_1057_out0 = v_G1_4365_out0;
assign v__2035_out0 = { v__5811_out0,v_S_1365_out0 };
assign v__2050_out0 = { v__5826_out0,v_S_1589_out0 };
assign v_CIN_9942_out0 = v_COUT_833_out0;
assign v_CIN_10166_out0 = v_COUT_1057_out0;
assign v_RD_6141_out0 = v_CIN_9942_out0;
assign v_RD_6605_out0 = v_CIN_10166_out0;
assign v_G1_7996_out0 = ((v_RD_6141_out0 && !v_RM_11581_out0) || (!v_RD_6141_out0) && v_RM_11581_out0);
assign v_G1_8460_out0 = ((v_RD_6605_out0 && !v_RM_12045_out0) || (!v_RD_6605_out0) && v_RM_12045_out0);
assign v_G2_12532_out0 = v_RD_6141_out0 && v_RM_11581_out0;
assign v_G2_12996_out0 = v_RD_6605_out0 && v_RM_12045_out0;
assign v_CARRY_5141_out0 = v_G2_12532_out0;
assign v_CARRY_5605_out0 = v_G2_12996_out0;
assign v_S_9142_out0 = v_G1_7996_out0;
assign v_S_9606_out0 = v_G1_8460_out0;
assign v_S_1353_out0 = v_S_9142_out0;
assign v_S_1577_out0 = v_S_9606_out0;
assign v_G1_4129_out0 = v_CARRY_5141_out0 || v_CARRY_5140_out0;
assign v_G1_4353_out0 = v_CARRY_5605_out0 || v_CARRY_5604_out0;
assign v_COUT_821_out0 = v_G1_4129_out0;
assign v_COUT_1045_out0 = v_G1_4353_out0;
assign v__2802_out0 = { v__2035_out0,v_S_1353_out0 };
assign v__2817_out0 = { v__2050_out0,v_S_1577_out0 };
assign v_CIN_9947_out0 = v_COUT_821_out0;
assign v_CIN_10171_out0 = v_COUT_1045_out0;
assign v_RD_6151_out0 = v_CIN_9947_out0;
assign v_RD_6615_out0 = v_CIN_10171_out0;
assign v_G1_8006_out0 = ((v_RD_6151_out0 && !v_RM_11591_out0) || (!v_RD_6151_out0) && v_RM_11591_out0);
assign v_G1_8470_out0 = ((v_RD_6615_out0 && !v_RM_12055_out0) || (!v_RD_6615_out0) && v_RM_12055_out0);
assign v_G2_12542_out0 = v_RD_6151_out0 && v_RM_11591_out0;
assign v_G2_13006_out0 = v_RD_6615_out0 && v_RM_12055_out0;
assign v_CARRY_5151_out0 = v_G2_12542_out0;
assign v_CARRY_5615_out0 = v_G2_13006_out0;
assign v_S_9152_out0 = v_G1_8006_out0;
assign v_S_9616_out0 = v_G1_8470_out0;
assign v_S_1358_out0 = v_S_9152_out0;
assign v_S_1582_out0 = v_S_9616_out0;
assign v_G1_4134_out0 = v_CARRY_5151_out0 || v_CARRY_5150_out0;
assign v_G1_4358_out0 = v_CARRY_5615_out0 || v_CARRY_5614_out0;
assign v_COUT_826_out0 = v_G1_4134_out0;
assign v_COUT_1050_out0 = v_G1_4358_out0;
assign v__1834_out0 = { v__2802_out0,v_S_1358_out0 };
assign v__1849_out0 = { v__2817_out0,v_S_1582_out0 };
assign v_CIN_9943_out0 = v_COUT_826_out0;
assign v_CIN_10167_out0 = v_COUT_1050_out0;
assign v_RD_6143_out0 = v_CIN_9943_out0;
assign v_RD_6607_out0 = v_CIN_10167_out0;
assign v_G1_7998_out0 = ((v_RD_6143_out0 && !v_RM_11583_out0) || (!v_RD_6143_out0) && v_RM_11583_out0);
assign v_G1_8462_out0 = ((v_RD_6607_out0 && !v_RM_12047_out0) || (!v_RD_6607_out0) && v_RM_12047_out0);
assign v_G2_12534_out0 = v_RD_6143_out0 && v_RM_11583_out0;
assign v_G2_12998_out0 = v_RD_6607_out0 && v_RM_12047_out0;
assign v_CARRY_5143_out0 = v_G2_12534_out0;
assign v_CARRY_5607_out0 = v_G2_12998_out0;
assign v_S_9144_out0 = v_G1_7998_out0;
assign v_S_9608_out0 = v_G1_8462_out0;
assign v_S_1354_out0 = v_S_9144_out0;
assign v_S_1578_out0 = v_S_9608_out0;
assign v_G1_4130_out0 = v_CARRY_5143_out0 || v_CARRY_5142_out0;
assign v_G1_4354_out0 = v_CARRY_5607_out0 || v_CARRY_5606_out0;
assign v_COUT_822_out0 = v_G1_4130_out0;
assign v_COUT_1046_out0 = v_G1_4354_out0;
assign v__4558_out0 = { v__1834_out0,v_S_1354_out0 };
assign v__4573_out0 = { v__1849_out0,v_S_1578_out0 };
assign v_RM_3491_out0 = v_COUT_822_out0;
assign v_RM_3715_out0 = v_COUT_1046_out0;
assign v_RM_11584_out0 = v_RM_3491_out0;
assign v_RM_12048_out0 = v_RM_3715_out0;
assign v_G1_7999_out0 = ((v_RD_6144_out0 && !v_RM_11584_out0) || (!v_RD_6144_out0) && v_RM_11584_out0);
assign v_G1_8463_out0 = ((v_RD_6608_out0 && !v_RM_12048_out0) || (!v_RD_6608_out0) && v_RM_12048_out0);
assign v_G2_12535_out0 = v_RD_6144_out0 && v_RM_11584_out0;
assign v_G2_12999_out0 = v_RD_6608_out0 && v_RM_12048_out0;
assign v_CARRY_5144_out0 = v_G2_12535_out0;
assign v_CARRY_5608_out0 = v_G2_12999_out0;
assign v_S_9145_out0 = v_G1_7999_out0;
assign v_S_9609_out0 = v_G1_8463_out0;
assign v_RM_11585_out0 = v_S_9145_out0;
assign v_RM_12049_out0 = v_S_9609_out0;
assign v_G1_8000_out0 = ((v_RD_6145_out0 && !v_RM_11585_out0) || (!v_RD_6145_out0) && v_RM_11585_out0);
assign v_G1_8464_out0 = ((v_RD_6609_out0 && !v_RM_12049_out0) || (!v_RD_6609_out0) && v_RM_12049_out0);
assign v_G2_12536_out0 = v_RD_6145_out0 && v_RM_11585_out0;
assign v_G2_13000_out0 = v_RD_6609_out0 && v_RM_12049_out0;
assign v_CARRY_5145_out0 = v_G2_12536_out0;
assign v_CARRY_5609_out0 = v_G2_13000_out0;
assign v_S_9146_out0 = v_G1_8000_out0;
assign v_S_9610_out0 = v_G1_8464_out0;
assign v_S_1355_out0 = v_S_9146_out0;
assign v_S_1579_out0 = v_S_9610_out0;
assign v_G1_4131_out0 = v_CARRY_5145_out0 || v_CARRY_5144_out0;
assign v_G1_4355_out0 = v_CARRY_5609_out0 || v_CARRY_5608_out0;
assign v_COUT_823_out0 = v_G1_4131_out0;
assign v_COUT_1047_out0 = v_G1_4355_out0;
assign v__10660_out0 = { v__4558_out0,v_S_1355_out0 };
assign v__10675_out0 = { v__4573_out0,v_S_1579_out0 };
assign v__10955_out0 = { v__10660_out0,v_COUT_823_out0 };
assign v__10970_out0 = { v__10675_out0,v_COUT_1047_out0 };
assign v_COUT_10925_out0 = v__10955_out0;
assign v_COUT_10940_out0 = v__10970_out0;
assign v_CIN_2369_out0 = v_COUT_10925_out0;
assign v_CIN_2384_out0 = v_COUT_10940_out0;
assign v__482_out0 = v_CIN_2369_out0[8:8];
assign v__497_out0 = v_CIN_2384_out0[8:8];
assign v__1787_out0 = v_CIN_2369_out0[6:6];
assign v__1802_out0 = v_CIN_2384_out0[6:6];
assign v__2169_out0 = v_CIN_2369_out0[3:3];
assign v__2184_out0 = v_CIN_2384_out0[3:3];
assign v__2208_out0 = v_CIN_2369_out0[15:15];
assign v__2222_out0 = v_CIN_2384_out0[15:15];
assign v__2516_out0 = v_CIN_2369_out0[0:0];
assign v__2531_out0 = v_CIN_2384_out0[0:0];
assign v__3065_out0 = v_CIN_2369_out0[9:9];
assign v__3080_out0 = v_CIN_2384_out0[9:9];
assign v__3099_out0 = v_CIN_2369_out0[2:2];
assign v__3114_out0 = v_CIN_2384_out0[2:2];
assign v__3153_out0 = v_CIN_2369_out0[7:7];
assign v__3168_out0 = v_CIN_2384_out0[7:7];
assign v__3837_out0 = v_CIN_2369_out0[1:1];
assign v__3852_out0 = v_CIN_2384_out0[1:1];
assign v__3875_out0 = v_CIN_2369_out0[10:10];
assign v__3890_out0 = v_CIN_2384_out0[10:10];
assign v__6814_out0 = v_CIN_2369_out0[11:11];
assign v__6829_out0 = v_CIN_2384_out0[11:11];
assign v__7658_out0 = v_CIN_2369_out0[12:12];
assign v__7673_out0 = v_CIN_2384_out0[12:12];
assign v__8713_out0 = v_CIN_2369_out0[13:13];
assign v__8728_out0 = v_CIN_2384_out0[13:13];
assign v__8783_out0 = v_CIN_2369_out0[14:14];
assign v__8798_out0 = v_CIN_2384_out0[14:14];
assign v__10733_out0 = v_CIN_2369_out0[5:5];
assign v__10748_out0 = v_CIN_2384_out0[5:5];
assign v__13462_out0 = v_CIN_2369_out0[4:4];
assign v__13477_out0 = v_CIN_2384_out0[4:4];
assign v_RM_3564_out0 = v__7658_out0;
assign v_RM_3565_out0 = v__8783_out0;
assign v_RM_3567_out0 = v__10733_out0;
assign v_RM_3568_out0 = v__13462_out0;
assign v_RM_3569_out0 = v__8713_out0;
assign v_RM_3570_out0 = v__3065_out0;
assign v_RM_3571_out0 = v__3875_out0;
assign v_RM_3572_out0 = v__3837_out0;
assign v_RM_3573_out0 = v__2169_out0;
assign v_RM_3574_out0 = v__1787_out0;
assign v_RM_3575_out0 = v__3153_out0;
assign v_RM_3576_out0 = v__6814_out0;
assign v_RM_3577_out0 = v__482_out0;
assign v_RM_3578_out0 = v__3099_out0;
assign v_RM_3788_out0 = v__7673_out0;
assign v_RM_3789_out0 = v__8798_out0;
assign v_RM_3791_out0 = v__10748_out0;
assign v_RM_3792_out0 = v__13477_out0;
assign v_RM_3793_out0 = v__8728_out0;
assign v_RM_3794_out0 = v__3080_out0;
assign v_RM_3795_out0 = v__3890_out0;
assign v_RM_3796_out0 = v__3852_out0;
assign v_RM_3797_out0 = v__2184_out0;
assign v_RM_3798_out0 = v__1802_out0;
assign v_RM_3799_out0 = v__3168_out0;
assign v_RM_3800_out0 = v__6829_out0;
assign v_RM_3801_out0 = v__497_out0;
assign v_RM_3802_out0 = v__3114_out0;
assign v_CIN_10019_out0 = v__2208_out0;
assign v_CIN_10243_out0 = v__2222_out0;
assign v_RM_11747_out0 = v__2516_out0;
assign v_RM_12211_out0 = v__2531_out0;
assign v_RD_6300_out0 = v_CIN_10019_out0;
assign v_RD_6764_out0 = v_CIN_10243_out0;
assign v_G1_8162_out0 = ((v_RD_6307_out0 && !v_RM_11747_out0) || (!v_RD_6307_out0) && v_RM_11747_out0);
assign v_G1_8626_out0 = ((v_RD_6771_out0 && !v_RM_12211_out0) || (!v_RD_6771_out0) && v_RM_12211_out0);
assign v_RM_11735_out0 = v_RM_3564_out0;
assign v_RM_11737_out0 = v_RM_3565_out0;
assign v_RM_11741_out0 = v_RM_3567_out0;
assign v_RM_11743_out0 = v_RM_3568_out0;
assign v_RM_11745_out0 = v_RM_3569_out0;
assign v_RM_11748_out0 = v_RM_3570_out0;
assign v_RM_11750_out0 = v_RM_3571_out0;
assign v_RM_11752_out0 = v_RM_3572_out0;
assign v_RM_11754_out0 = v_RM_3573_out0;
assign v_RM_11756_out0 = v_RM_3574_out0;
assign v_RM_11758_out0 = v_RM_3575_out0;
assign v_RM_11760_out0 = v_RM_3576_out0;
assign v_RM_11762_out0 = v_RM_3577_out0;
assign v_RM_11764_out0 = v_RM_3578_out0;
assign v_RM_12199_out0 = v_RM_3788_out0;
assign v_RM_12201_out0 = v_RM_3789_out0;
assign v_RM_12205_out0 = v_RM_3791_out0;
assign v_RM_12207_out0 = v_RM_3792_out0;
assign v_RM_12209_out0 = v_RM_3793_out0;
assign v_RM_12212_out0 = v_RM_3794_out0;
assign v_RM_12214_out0 = v_RM_3795_out0;
assign v_RM_12216_out0 = v_RM_3796_out0;
assign v_RM_12218_out0 = v_RM_3797_out0;
assign v_RM_12220_out0 = v_RM_3798_out0;
assign v_RM_12222_out0 = v_RM_3799_out0;
assign v_RM_12224_out0 = v_RM_3800_out0;
assign v_RM_12226_out0 = v_RM_3801_out0;
assign v_RM_12228_out0 = v_RM_3802_out0;
assign v_G2_12698_out0 = v_RD_6307_out0 && v_RM_11747_out0;
assign v_G2_13162_out0 = v_RD_6771_out0 && v_RM_12211_out0;
assign v_CARRY_5307_out0 = v_G2_12698_out0;
assign v_CARRY_5771_out0 = v_G2_13162_out0;
assign v_G1_8150_out0 = ((v_RD_6295_out0 && !v_RM_11735_out0) || (!v_RD_6295_out0) && v_RM_11735_out0);
assign v_G1_8152_out0 = ((v_RD_6297_out0 && !v_RM_11737_out0) || (!v_RD_6297_out0) && v_RM_11737_out0);
assign v_G1_8156_out0 = ((v_RD_6301_out0 && !v_RM_11741_out0) || (!v_RD_6301_out0) && v_RM_11741_out0);
assign v_G1_8158_out0 = ((v_RD_6303_out0 && !v_RM_11743_out0) || (!v_RD_6303_out0) && v_RM_11743_out0);
assign v_G1_8160_out0 = ((v_RD_6305_out0 && !v_RM_11745_out0) || (!v_RD_6305_out0) && v_RM_11745_out0);
assign v_G1_8163_out0 = ((v_RD_6308_out0 && !v_RM_11748_out0) || (!v_RD_6308_out0) && v_RM_11748_out0);
assign v_G1_8165_out0 = ((v_RD_6310_out0 && !v_RM_11750_out0) || (!v_RD_6310_out0) && v_RM_11750_out0);
assign v_G1_8167_out0 = ((v_RD_6312_out0 && !v_RM_11752_out0) || (!v_RD_6312_out0) && v_RM_11752_out0);
assign v_G1_8169_out0 = ((v_RD_6314_out0 && !v_RM_11754_out0) || (!v_RD_6314_out0) && v_RM_11754_out0);
assign v_G1_8171_out0 = ((v_RD_6316_out0 && !v_RM_11756_out0) || (!v_RD_6316_out0) && v_RM_11756_out0);
assign v_G1_8173_out0 = ((v_RD_6318_out0 && !v_RM_11758_out0) || (!v_RD_6318_out0) && v_RM_11758_out0);
assign v_G1_8175_out0 = ((v_RD_6320_out0 && !v_RM_11760_out0) || (!v_RD_6320_out0) && v_RM_11760_out0);
assign v_G1_8177_out0 = ((v_RD_6322_out0 && !v_RM_11762_out0) || (!v_RD_6322_out0) && v_RM_11762_out0);
assign v_G1_8179_out0 = ((v_RD_6324_out0 && !v_RM_11764_out0) || (!v_RD_6324_out0) && v_RM_11764_out0);
assign v_G1_8614_out0 = ((v_RD_6759_out0 && !v_RM_12199_out0) || (!v_RD_6759_out0) && v_RM_12199_out0);
assign v_G1_8616_out0 = ((v_RD_6761_out0 && !v_RM_12201_out0) || (!v_RD_6761_out0) && v_RM_12201_out0);
assign v_G1_8620_out0 = ((v_RD_6765_out0 && !v_RM_12205_out0) || (!v_RD_6765_out0) && v_RM_12205_out0);
assign v_G1_8622_out0 = ((v_RD_6767_out0 && !v_RM_12207_out0) || (!v_RD_6767_out0) && v_RM_12207_out0);
assign v_G1_8624_out0 = ((v_RD_6769_out0 && !v_RM_12209_out0) || (!v_RD_6769_out0) && v_RM_12209_out0);
assign v_G1_8627_out0 = ((v_RD_6772_out0 && !v_RM_12212_out0) || (!v_RD_6772_out0) && v_RM_12212_out0);
assign v_G1_8629_out0 = ((v_RD_6774_out0 && !v_RM_12214_out0) || (!v_RD_6774_out0) && v_RM_12214_out0);
assign v_G1_8631_out0 = ((v_RD_6776_out0 && !v_RM_12216_out0) || (!v_RD_6776_out0) && v_RM_12216_out0);
assign v_G1_8633_out0 = ((v_RD_6778_out0 && !v_RM_12218_out0) || (!v_RD_6778_out0) && v_RM_12218_out0);
assign v_G1_8635_out0 = ((v_RD_6780_out0 && !v_RM_12220_out0) || (!v_RD_6780_out0) && v_RM_12220_out0);
assign v_G1_8637_out0 = ((v_RD_6782_out0 && !v_RM_12222_out0) || (!v_RD_6782_out0) && v_RM_12222_out0);
assign v_G1_8639_out0 = ((v_RD_6784_out0 && !v_RM_12224_out0) || (!v_RD_6784_out0) && v_RM_12224_out0);
assign v_G1_8641_out0 = ((v_RD_6786_out0 && !v_RM_12226_out0) || (!v_RD_6786_out0) && v_RM_12226_out0);
assign v_G1_8643_out0 = ((v_RD_6788_out0 && !v_RM_12228_out0) || (!v_RD_6788_out0) && v_RM_12228_out0);
assign v_S_9308_out0 = v_G1_8162_out0;
assign v_S_9772_out0 = v_G1_8626_out0;
assign v_G2_12686_out0 = v_RD_6295_out0 && v_RM_11735_out0;
assign v_G2_12688_out0 = v_RD_6297_out0 && v_RM_11737_out0;
assign v_G2_12692_out0 = v_RD_6301_out0 && v_RM_11741_out0;
assign v_G2_12694_out0 = v_RD_6303_out0 && v_RM_11743_out0;
assign v_G2_12696_out0 = v_RD_6305_out0 && v_RM_11745_out0;
assign v_G2_12699_out0 = v_RD_6308_out0 && v_RM_11748_out0;
assign v_G2_12701_out0 = v_RD_6310_out0 && v_RM_11750_out0;
assign v_G2_12703_out0 = v_RD_6312_out0 && v_RM_11752_out0;
assign v_G2_12705_out0 = v_RD_6314_out0 && v_RM_11754_out0;
assign v_G2_12707_out0 = v_RD_6316_out0 && v_RM_11756_out0;
assign v_G2_12709_out0 = v_RD_6318_out0 && v_RM_11758_out0;
assign v_G2_12711_out0 = v_RD_6320_out0 && v_RM_11760_out0;
assign v_G2_12713_out0 = v_RD_6322_out0 && v_RM_11762_out0;
assign v_G2_12715_out0 = v_RD_6324_out0 && v_RM_11764_out0;
assign v_G2_13150_out0 = v_RD_6759_out0 && v_RM_12199_out0;
assign v_G2_13152_out0 = v_RD_6761_out0 && v_RM_12201_out0;
assign v_G2_13156_out0 = v_RD_6765_out0 && v_RM_12205_out0;
assign v_G2_13158_out0 = v_RD_6767_out0 && v_RM_12207_out0;
assign v_G2_13160_out0 = v_RD_6769_out0 && v_RM_12209_out0;
assign v_G2_13163_out0 = v_RD_6772_out0 && v_RM_12212_out0;
assign v_G2_13165_out0 = v_RD_6774_out0 && v_RM_12214_out0;
assign v_G2_13167_out0 = v_RD_6776_out0 && v_RM_12216_out0;
assign v_G2_13169_out0 = v_RD_6778_out0 && v_RM_12218_out0;
assign v_G2_13171_out0 = v_RD_6780_out0 && v_RM_12220_out0;
assign v_G2_13173_out0 = v_RD_6782_out0 && v_RM_12222_out0;
assign v_G2_13175_out0 = v_RD_6784_out0 && v_RM_12224_out0;
assign v_G2_13177_out0 = v_RD_6786_out0 && v_RM_12226_out0;
assign v_G2_13179_out0 = v_RD_6788_out0 && v_RM_12228_out0;
assign v_S_4679_out0 = v_S_9308_out0;
assign v_S_4694_out0 = v_S_9772_out0;
assign v_CARRY_5295_out0 = v_G2_12686_out0;
assign v_CARRY_5297_out0 = v_G2_12688_out0;
assign v_CARRY_5301_out0 = v_G2_12692_out0;
assign v_CARRY_5303_out0 = v_G2_12694_out0;
assign v_CARRY_5305_out0 = v_G2_12696_out0;
assign v_CARRY_5308_out0 = v_G2_12699_out0;
assign v_CARRY_5310_out0 = v_G2_12701_out0;
assign v_CARRY_5312_out0 = v_G2_12703_out0;
assign v_CARRY_5314_out0 = v_G2_12705_out0;
assign v_CARRY_5316_out0 = v_G2_12707_out0;
assign v_CARRY_5318_out0 = v_G2_12709_out0;
assign v_CARRY_5320_out0 = v_G2_12711_out0;
assign v_CARRY_5322_out0 = v_G2_12713_out0;
assign v_CARRY_5324_out0 = v_G2_12715_out0;
assign v_CARRY_5759_out0 = v_G2_13150_out0;
assign v_CARRY_5761_out0 = v_G2_13152_out0;
assign v_CARRY_5765_out0 = v_G2_13156_out0;
assign v_CARRY_5767_out0 = v_G2_13158_out0;
assign v_CARRY_5769_out0 = v_G2_13160_out0;
assign v_CARRY_5772_out0 = v_G2_13163_out0;
assign v_CARRY_5774_out0 = v_G2_13165_out0;
assign v_CARRY_5776_out0 = v_G2_13167_out0;
assign v_CARRY_5778_out0 = v_G2_13169_out0;
assign v_CARRY_5780_out0 = v_G2_13171_out0;
assign v_CARRY_5782_out0 = v_G2_13173_out0;
assign v_CARRY_5784_out0 = v_G2_13175_out0;
assign v_CARRY_5786_out0 = v_G2_13177_out0;
assign v_CARRY_5788_out0 = v_G2_13179_out0;
assign v_S_9296_out0 = v_G1_8150_out0;
assign v_S_9298_out0 = v_G1_8152_out0;
assign v_S_9302_out0 = v_G1_8156_out0;
assign v_S_9304_out0 = v_G1_8158_out0;
assign v_S_9306_out0 = v_G1_8160_out0;
assign v_S_9309_out0 = v_G1_8163_out0;
assign v_S_9311_out0 = v_G1_8165_out0;
assign v_S_9313_out0 = v_G1_8167_out0;
assign v_S_9315_out0 = v_G1_8169_out0;
assign v_S_9317_out0 = v_G1_8171_out0;
assign v_S_9319_out0 = v_G1_8173_out0;
assign v_S_9321_out0 = v_G1_8175_out0;
assign v_S_9323_out0 = v_G1_8177_out0;
assign v_S_9325_out0 = v_G1_8179_out0;
assign v_S_9760_out0 = v_G1_8614_out0;
assign v_S_9762_out0 = v_G1_8616_out0;
assign v_S_9766_out0 = v_G1_8620_out0;
assign v_S_9768_out0 = v_G1_8622_out0;
assign v_S_9770_out0 = v_G1_8624_out0;
assign v_S_9773_out0 = v_G1_8627_out0;
assign v_S_9775_out0 = v_G1_8629_out0;
assign v_S_9777_out0 = v_G1_8631_out0;
assign v_S_9779_out0 = v_G1_8633_out0;
assign v_S_9781_out0 = v_G1_8635_out0;
assign v_S_9783_out0 = v_G1_8637_out0;
assign v_S_9785_out0 = v_G1_8639_out0;
assign v_S_9787_out0 = v_G1_8641_out0;
assign v_S_9789_out0 = v_G1_8643_out0;
assign v_CIN_10025_out0 = v_CARRY_5307_out0;
assign v_CIN_10249_out0 = v_CARRY_5771_out0;
assign v_RD_6313_out0 = v_CIN_10025_out0;
assign v_RD_6777_out0 = v_CIN_10249_out0;
assign v__10775_out0 = { v__43_out0,v_S_4679_out0 };
assign v__10776_out0 = { v__44_out0,v_S_4694_out0 };
assign v_RM_11736_out0 = v_S_9296_out0;
assign v_RM_11738_out0 = v_S_9298_out0;
assign v_RM_11742_out0 = v_S_9302_out0;
assign v_RM_11744_out0 = v_S_9304_out0;
assign v_RM_11746_out0 = v_S_9306_out0;
assign v_RM_11749_out0 = v_S_9309_out0;
assign v_RM_11751_out0 = v_S_9311_out0;
assign v_RM_11753_out0 = v_S_9313_out0;
assign v_RM_11755_out0 = v_S_9315_out0;
assign v_RM_11757_out0 = v_S_9317_out0;
assign v_RM_11759_out0 = v_S_9319_out0;
assign v_RM_11761_out0 = v_S_9321_out0;
assign v_RM_11763_out0 = v_S_9323_out0;
assign v_RM_11765_out0 = v_S_9325_out0;
assign v_RM_12200_out0 = v_S_9760_out0;
assign v_RM_12202_out0 = v_S_9762_out0;
assign v_RM_12206_out0 = v_S_9766_out0;
assign v_RM_12208_out0 = v_S_9768_out0;
assign v_RM_12210_out0 = v_S_9770_out0;
assign v_RM_12213_out0 = v_S_9773_out0;
assign v_RM_12215_out0 = v_S_9775_out0;
assign v_RM_12217_out0 = v_S_9777_out0;
assign v_RM_12219_out0 = v_S_9779_out0;
assign v_RM_12221_out0 = v_S_9781_out0;
assign v_RM_12223_out0 = v_S_9783_out0;
assign v_RM_12225_out0 = v_S_9785_out0;
assign v_RM_12227_out0 = v_S_9787_out0;
assign v_RM_12229_out0 = v_S_9789_out0;
assign v_G1_8168_out0 = ((v_RD_6313_out0 && !v_RM_11753_out0) || (!v_RD_6313_out0) && v_RM_11753_out0);
assign v_G1_8632_out0 = ((v_RD_6777_out0 && !v_RM_12217_out0) || (!v_RD_6777_out0) && v_RM_12217_out0);
assign v_G2_12704_out0 = v_RD_6313_out0 && v_RM_11753_out0;
assign v_G2_13168_out0 = v_RD_6777_out0 && v_RM_12217_out0;
assign v_CARRY_5313_out0 = v_G2_12704_out0;
assign v_CARRY_5777_out0 = v_G2_13168_out0;
assign v_S_9314_out0 = v_G1_8168_out0;
assign v_S_9778_out0 = v_G1_8632_out0;
assign v_S_1436_out0 = v_S_9314_out0;
assign v_S_1660_out0 = v_S_9778_out0;
assign v_G1_4212_out0 = v_CARRY_5313_out0 || v_CARRY_5312_out0;
assign v_G1_4436_out0 = v_CARRY_5777_out0 || v_CARRY_5776_out0;
assign v_COUT_904_out0 = v_G1_4212_out0;
assign v_COUT_1128_out0 = v_G1_4436_out0;
assign v_CIN_10031_out0 = v_COUT_904_out0;
assign v_CIN_10255_out0 = v_COUT_1128_out0;
assign v_RD_6325_out0 = v_CIN_10031_out0;
assign v_RD_6789_out0 = v_CIN_10255_out0;
assign v_G1_8180_out0 = ((v_RD_6325_out0 && !v_RM_11765_out0) || (!v_RD_6325_out0) && v_RM_11765_out0);
assign v_G1_8644_out0 = ((v_RD_6789_out0 && !v_RM_12229_out0) || (!v_RD_6789_out0) && v_RM_12229_out0);
assign v_G2_12716_out0 = v_RD_6325_out0 && v_RM_11765_out0;
assign v_G2_13180_out0 = v_RD_6789_out0 && v_RM_12229_out0;
assign v_CARRY_5325_out0 = v_G2_12716_out0;
assign v_CARRY_5789_out0 = v_G2_13180_out0;
assign v_S_9326_out0 = v_G1_8180_out0;
assign v_S_9790_out0 = v_G1_8644_out0;
assign v_S_1442_out0 = v_S_9326_out0;
assign v_S_1666_out0 = v_S_9790_out0;
assign v_G1_4218_out0 = v_CARRY_5325_out0 || v_CARRY_5324_out0;
assign v_G1_4442_out0 = v_CARRY_5789_out0 || v_CARRY_5788_out0;
assign v_COUT_910_out0 = v_G1_4218_out0;
assign v_COUT_1134_out0 = v_G1_4442_out0;
assign v__4796_out0 = { v_S_1436_out0,v_S_1442_out0 };
assign v__4811_out0 = { v_S_1660_out0,v_S_1666_out0 };
assign v_CIN_10026_out0 = v_COUT_910_out0;
assign v_CIN_10250_out0 = v_COUT_1134_out0;
assign v_RD_6315_out0 = v_CIN_10026_out0;
assign v_RD_6779_out0 = v_CIN_10250_out0;
assign v_G1_8170_out0 = ((v_RD_6315_out0 && !v_RM_11755_out0) || (!v_RD_6315_out0) && v_RM_11755_out0);
assign v_G1_8634_out0 = ((v_RD_6779_out0 && !v_RM_12219_out0) || (!v_RD_6779_out0) && v_RM_12219_out0);
assign v_G2_12706_out0 = v_RD_6315_out0 && v_RM_11755_out0;
assign v_G2_13170_out0 = v_RD_6779_out0 && v_RM_12219_out0;
assign v_CARRY_5315_out0 = v_G2_12706_out0;
assign v_CARRY_5779_out0 = v_G2_13170_out0;
assign v_S_9316_out0 = v_G1_8170_out0;
assign v_S_9780_out0 = v_G1_8634_out0;
assign v_S_1437_out0 = v_S_9316_out0;
assign v_S_1661_out0 = v_S_9780_out0;
assign v_G1_4213_out0 = v_CARRY_5315_out0 || v_CARRY_5314_out0;
assign v_G1_4437_out0 = v_CARRY_5779_out0 || v_CARRY_5778_out0;
assign v_COUT_905_out0 = v_G1_4213_out0;
assign v_COUT_1129_out0 = v_G1_4437_out0;
assign v__2566_out0 = { v__4796_out0,v_S_1437_out0 };
assign v__2581_out0 = { v__4811_out0,v_S_1661_out0 };
assign v_CIN_10021_out0 = v_COUT_905_out0;
assign v_CIN_10245_out0 = v_COUT_1129_out0;
assign v_RD_6304_out0 = v_CIN_10021_out0;
assign v_RD_6768_out0 = v_CIN_10245_out0;
assign v_G1_8159_out0 = ((v_RD_6304_out0 && !v_RM_11744_out0) || (!v_RD_6304_out0) && v_RM_11744_out0);
assign v_G1_8623_out0 = ((v_RD_6768_out0 && !v_RM_12208_out0) || (!v_RD_6768_out0) && v_RM_12208_out0);
assign v_G2_12695_out0 = v_RD_6304_out0 && v_RM_11744_out0;
assign v_G2_13159_out0 = v_RD_6768_out0 && v_RM_12208_out0;
assign v_CARRY_5304_out0 = v_G2_12695_out0;
assign v_CARRY_5768_out0 = v_G2_13159_out0;
assign v_S_9305_out0 = v_G1_8159_out0;
assign v_S_9769_out0 = v_G1_8623_out0;
assign v_S_1432_out0 = v_S_9305_out0;
assign v_S_1656_out0 = v_S_9769_out0;
assign v_G1_4208_out0 = v_CARRY_5304_out0 || v_CARRY_5303_out0;
assign v_G1_4432_out0 = v_CARRY_5768_out0 || v_CARRY_5767_out0;
assign v_COUT_900_out0 = v_G1_4208_out0;
assign v_COUT_1124_out0 = v_G1_4432_out0;
assign v__7046_out0 = { v__2566_out0,v_S_1432_out0 };
assign v__7061_out0 = { v__2581_out0,v_S_1656_out0 };
assign v_CIN_10020_out0 = v_COUT_900_out0;
assign v_CIN_10244_out0 = v_COUT_1124_out0;
assign v_RD_6302_out0 = v_CIN_10020_out0;
assign v_RD_6766_out0 = v_CIN_10244_out0;
assign v_G1_8157_out0 = ((v_RD_6302_out0 && !v_RM_11742_out0) || (!v_RD_6302_out0) && v_RM_11742_out0);
assign v_G1_8621_out0 = ((v_RD_6766_out0 && !v_RM_12206_out0) || (!v_RD_6766_out0) && v_RM_12206_out0);
assign v_G2_12693_out0 = v_RD_6302_out0 && v_RM_11742_out0;
assign v_G2_13157_out0 = v_RD_6766_out0 && v_RM_12206_out0;
assign v_CARRY_5302_out0 = v_G2_12693_out0;
assign v_CARRY_5766_out0 = v_G2_13157_out0;
assign v_S_9303_out0 = v_G1_8157_out0;
assign v_S_9767_out0 = v_G1_8621_out0;
assign v_S_1431_out0 = v_S_9303_out0;
assign v_S_1655_out0 = v_S_9767_out0;
assign v_G1_4207_out0 = v_CARRY_5302_out0 || v_CARRY_5301_out0;
assign v_G1_4431_out0 = v_CARRY_5766_out0 || v_CARRY_5765_out0;
assign v_COUT_899_out0 = v_G1_4207_out0;
assign v_COUT_1123_out0 = v_G1_4431_out0;
assign v__13532_out0 = { v__7046_out0,v_S_1431_out0 };
assign v__13547_out0 = { v__7061_out0,v_S_1655_out0 };
assign v_CIN_10027_out0 = v_COUT_899_out0;
assign v_CIN_10251_out0 = v_COUT_1123_out0;
assign v_RD_6317_out0 = v_CIN_10027_out0;
assign v_RD_6781_out0 = v_CIN_10251_out0;
assign v_G1_8172_out0 = ((v_RD_6317_out0 && !v_RM_11757_out0) || (!v_RD_6317_out0) && v_RM_11757_out0);
assign v_G1_8636_out0 = ((v_RD_6781_out0 && !v_RM_12221_out0) || (!v_RD_6781_out0) && v_RM_12221_out0);
assign v_G2_12708_out0 = v_RD_6317_out0 && v_RM_11757_out0;
assign v_G2_13172_out0 = v_RD_6781_out0 && v_RM_12221_out0;
assign v_CARRY_5317_out0 = v_G2_12708_out0;
assign v_CARRY_5781_out0 = v_G2_13172_out0;
assign v_S_9318_out0 = v_G1_8172_out0;
assign v_S_9782_out0 = v_G1_8636_out0;
assign v_S_1438_out0 = v_S_9318_out0;
assign v_S_1662_out0 = v_S_9782_out0;
assign v_G1_4214_out0 = v_CARRY_5317_out0 || v_CARRY_5316_out0;
assign v_G1_4438_out0 = v_CARRY_5781_out0 || v_CARRY_5780_out0;
assign v_COUT_906_out0 = v_G1_4214_out0;
assign v_COUT_1130_out0 = v_G1_4438_out0;
assign v__3325_out0 = { v__13532_out0,v_S_1438_out0 };
assign v__3340_out0 = { v__13547_out0,v_S_1662_out0 };
assign v_CIN_10028_out0 = v_COUT_906_out0;
assign v_CIN_10252_out0 = v_COUT_1130_out0;
assign v_RD_6319_out0 = v_CIN_10028_out0;
assign v_RD_6783_out0 = v_CIN_10252_out0;
assign v_G1_8174_out0 = ((v_RD_6319_out0 && !v_RM_11759_out0) || (!v_RD_6319_out0) && v_RM_11759_out0);
assign v_G1_8638_out0 = ((v_RD_6783_out0 && !v_RM_12223_out0) || (!v_RD_6783_out0) && v_RM_12223_out0);
assign v_G2_12710_out0 = v_RD_6319_out0 && v_RM_11759_out0;
assign v_G2_13174_out0 = v_RD_6783_out0 && v_RM_12223_out0;
assign v_CARRY_5319_out0 = v_G2_12710_out0;
assign v_CARRY_5783_out0 = v_G2_13174_out0;
assign v_S_9320_out0 = v_G1_8174_out0;
assign v_S_9784_out0 = v_G1_8638_out0;
assign v_S_1439_out0 = v_S_9320_out0;
assign v_S_1663_out0 = v_S_9784_out0;
assign v_G1_4215_out0 = v_CARRY_5319_out0 || v_CARRY_5318_out0;
assign v_G1_4439_out0 = v_CARRY_5783_out0 || v_CARRY_5782_out0;
assign v_COUT_907_out0 = v_G1_4215_out0;
assign v_COUT_1131_out0 = v_G1_4439_out0;
assign v__7161_out0 = { v__3325_out0,v_S_1439_out0 };
assign v__7176_out0 = { v__3340_out0,v_S_1663_out0 };
assign v_CIN_10030_out0 = v_COUT_907_out0;
assign v_CIN_10254_out0 = v_COUT_1131_out0;
assign v_RD_6323_out0 = v_CIN_10030_out0;
assign v_RD_6787_out0 = v_CIN_10254_out0;
assign v_G1_8178_out0 = ((v_RD_6323_out0 && !v_RM_11763_out0) || (!v_RD_6323_out0) && v_RM_11763_out0);
assign v_G1_8642_out0 = ((v_RD_6787_out0 && !v_RM_12227_out0) || (!v_RD_6787_out0) && v_RM_12227_out0);
assign v_G2_12714_out0 = v_RD_6323_out0 && v_RM_11763_out0;
assign v_G2_13178_out0 = v_RD_6787_out0 && v_RM_12227_out0;
assign v_CARRY_5323_out0 = v_G2_12714_out0;
assign v_CARRY_5787_out0 = v_G2_13178_out0;
assign v_S_9324_out0 = v_G1_8178_out0;
assign v_S_9788_out0 = v_G1_8642_out0;
assign v_S_1441_out0 = v_S_9324_out0;
assign v_S_1665_out0 = v_S_9788_out0;
assign v_G1_4217_out0 = v_CARRY_5323_out0 || v_CARRY_5322_out0;
assign v_G1_4441_out0 = v_CARRY_5787_out0 || v_CARRY_5786_out0;
assign v_COUT_909_out0 = v_G1_4217_out0;
assign v_COUT_1133_out0 = v_G1_4441_out0;
assign v__4763_out0 = { v__7161_out0,v_S_1441_out0 };
assign v__4778_out0 = { v__7176_out0,v_S_1665_out0 };
assign v_CIN_10023_out0 = v_COUT_909_out0;
assign v_CIN_10247_out0 = v_COUT_1133_out0;
assign v_RD_6309_out0 = v_CIN_10023_out0;
assign v_RD_6773_out0 = v_CIN_10247_out0;
assign v_G1_8164_out0 = ((v_RD_6309_out0 && !v_RM_11749_out0) || (!v_RD_6309_out0) && v_RM_11749_out0);
assign v_G1_8628_out0 = ((v_RD_6773_out0 && !v_RM_12213_out0) || (!v_RD_6773_out0) && v_RM_12213_out0);
assign v_G2_12700_out0 = v_RD_6309_out0 && v_RM_11749_out0;
assign v_G2_13164_out0 = v_RD_6773_out0 && v_RM_12213_out0;
assign v_CARRY_5309_out0 = v_G2_12700_out0;
assign v_CARRY_5773_out0 = v_G2_13164_out0;
assign v_S_9310_out0 = v_G1_8164_out0;
assign v_S_9774_out0 = v_G1_8628_out0;
assign v_S_1434_out0 = v_S_9310_out0;
assign v_S_1658_out0 = v_S_9774_out0;
assign v_G1_4210_out0 = v_CARRY_5309_out0 || v_CARRY_5308_out0;
assign v_G1_4434_out0 = v_CARRY_5773_out0 || v_CARRY_5772_out0;
assign v_COUT_902_out0 = v_G1_4210_out0;
assign v_COUT_1126_out0 = v_G1_4434_out0;
assign v__6940_out0 = { v__4763_out0,v_S_1434_out0 };
assign v__6955_out0 = { v__4778_out0,v_S_1658_out0 };
assign v_CIN_10024_out0 = v_COUT_902_out0;
assign v_CIN_10248_out0 = v_COUT_1126_out0;
assign v_RD_6311_out0 = v_CIN_10024_out0;
assign v_RD_6775_out0 = v_CIN_10248_out0;
assign v_G1_8166_out0 = ((v_RD_6311_out0 && !v_RM_11751_out0) || (!v_RD_6311_out0) && v_RM_11751_out0);
assign v_G1_8630_out0 = ((v_RD_6775_out0 && !v_RM_12215_out0) || (!v_RD_6775_out0) && v_RM_12215_out0);
assign v_G2_12702_out0 = v_RD_6311_out0 && v_RM_11751_out0;
assign v_G2_13166_out0 = v_RD_6775_out0 && v_RM_12215_out0;
assign v_CARRY_5311_out0 = v_G2_12702_out0;
assign v_CARRY_5775_out0 = v_G2_13166_out0;
assign v_S_9312_out0 = v_G1_8166_out0;
assign v_S_9776_out0 = v_G1_8630_out0;
assign v_S_1435_out0 = v_S_9312_out0;
assign v_S_1659_out0 = v_S_9776_out0;
assign v_G1_4211_out0 = v_CARRY_5311_out0 || v_CARRY_5310_out0;
assign v_G1_4435_out0 = v_CARRY_5775_out0 || v_CARRY_5774_out0;
assign v_COUT_903_out0 = v_G1_4211_out0;
assign v_COUT_1127_out0 = v_G1_4435_out0;
assign v__5816_out0 = { v__6940_out0,v_S_1435_out0 };
assign v__5831_out0 = { v__6955_out0,v_S_1659_out0 };
assign v_CIN_10029_out0 = v_COUT_903_out0;
assign v_CIN_10253_out0 = v_COUT_1127_out0;
assign v_RD_6321_out0 = v_CIN_10029_out0;
assign v_RD_6785_out0 = v_CIN_10253_out0;
assign v_G1_8176_out0 = ((v_RD_6321_out0 && !v_RM_11761_out0) || (!v_RD_6321_out0) && v_RM_11761_out0);
assign v_G1_8640_out0 = ((v_RD_6785_out0 && !v_RM_12225_out0) || (!v_RD_6785_out0) && v_RM_12225_out0);
assign v_G2_12712_out0 = v_RD_6321_out0 && v_RM_11761_out0;
assign v_G2_13176_out0 = v_RD_6785_out0 && v_RM_12225_out0;
assign v_CARRY_5321_out0 = v_G2_12712_out0;
assign v_CARRY_5785_out0 = v_G2_13176_out0;
assign v_S_9322_out0 = v_G1_8176_out0;
assign v_S_9786_out0 = v_G1_8640_out0;
assign v_S_1440_out0 = v_S_9322_out0;
assign v_S_1664_out0 = v_S_9786_out0;
assign v_G1_4216_out0 = v_CARRY_5321_out0 || v_CARRY_5320_out0;
assign v_G1_4440_out0 = v_CARRY_5785_out0 || v_CARRY_5784_out0;
assign v_COUT_908_out0 = v_G1_4216_out0;
assign v_COUT_1132_out0 = v_G1_4440_out0;
assign v__2040_out0 = { v__5816_out0,v_S_1440_out0 };
assign v__2055_out0 = { v__5831_out0,v_S_1664_out0 };
assign v_CIN_10017_out0 = v_COUT_908_out0;
assign v_CIN_10241_out0 = v_COUT_1132_out0;
assign v_RD_6296_out0 = v_CIN_10017_out0;
assign v_RD_6760_out0 = v_CIN_10241_out0;
assign v_G1_8151_out0 = ((v_RD_6296_out0 && !v_RM_11736_out0) || (!v_RD_6296_out0) && v_RM_11736_out0);
assign v_G1_8615_out0 = ((v_RD_6760_out0 && !v_RM_12200_out0) || (!v_RD_6760_out0) && v_RM_12200_out0);
assign v_G2_12687_out0 = v_RD_6296_out0 && v_RM_11736_out0;
assign v_G2_13151_out0 = v_RD_6760_out0 && v_RM_12200_out0;
assign v_CARRY_5296_out0 = v_G2_12687_out0;
assign v_CARRY_5760_out0 = v_G2_13151_out0;
assign v_S_9297_out0 = v_G1_8151_out0;
assign v_S_9761_out0 = v_G1_8615_out0;
assign v_S_1428_out0 = v_S_9297_out0;
assign v_S_1652_out0 = v_S_9761_out0;
assign v_G1_4204_out0 = v_CARRY_5296_out0 || v_CARRY_5295_out0;
assign v_G1_4428_out0 = v_CARRY_5760_out0 || v_CARRY_5759_out0;
assign v_COUT_896_out0 = v_G1_4204_out0;
assign v_COUT_1120_out0 = v_G1_4428_out0;
assign v__2807_out0 = { v__2040_out0,v_S_1428_out0 };
assign v__2822_out0 = { v__2055_out0,v_S_1652_out0 };
assign v_CIN_10022_out0 = v_COUT_896_out0;
assign v_CIN_10246_out0 = v_COUT_1120_out0;
assign v_RD_6306_out0 = v_CIN_10022_out0;
assign v_RD_6770_out0 = v_CIN_10246_out0;
assign v_G1_8161_out0 = ((v_RD_6306_out0 && !v_RM_11746_out0) || (!v_RD_6306_out0) && v_RM_11746_out0);
assign v_G1_8625_out0 = ((v_RD_6770_out0 && !v_RM_12210_out0) || (!v_RD_6770_out0) && v_RM_12210_out0);
assign v_G2_12697_out0 = v_RD_6306_out0 && v_RM_11746_out0;
assign v_G2_13161_out0 = v_RD_6770_out0 && v_RM_12210_out0;
assign v_CARRY_5306_out0 = v_G2_12697_out0;
assign v_CARRY_5770_out0 = v_G2_13161_out0;
assign v_S_9307_out0 = v_G1_8161_out0;
assign v_S_9771_out0 = v_G1_8625_out0;
assign v_S_1433_out0 = v_S_9307_out0;
assign v_S_1657_out0 = v_S_9771_out0;
assign v_G1_4209_out0 = v_CARRY_5306_out0 || v_CARRY_5305_out0;
assign v_G1_4433_out0 = v_CARRY_5770_out0 || v_CARRY_5769_out0;
assign v_COUT_901_out0 = v_G1_4209_out0;
assign v_COUT_1125_out0 = v_G1_4433_out0;
assign v__1839_out0 = { v__2807_out0,v_S_1433_out0 };
assign v__1854_out0 = { v__2822_out0,v_S_1657_out0 };
assign v_CIN_10018_out0 = v_COUT_901_out0;
assign v_CIN_10242_out0 = v_COUT_1125_out0;
assign v_RD_6298_out0 = v_CIN_10018_out0;
assign v_RD_6762_out0 = v_CIN_10242_out0;
assign v_G1_8153_out0 = ((v_RD_6298_out0 && !v_RM_11738_out0) || (!v_RD_6298_out0) && v_RM_11738_out0);
assign v_G1_8617_out0 = ((v_RD_6762_out0 && !v_RM_12202_out0) || (!v_RD_6762_out0) && v_RM_12202_out0);
assign v_G2_12689_out0 = v_RD_6298_out0 && v_RM_11738_out0;
assign v_G2_13153_out0 = v_RD_6762_out0 && v_RM_12202_out0;
assign v_CARRY_5298_out0 = v_G2_12689_out0;
assign v_CARRY_5762_out0 = v_G2_13153_out0;
assign v_S_9299_out0 = v_G1_8153_out0;
assign v_S_9763_out0 = v_G1_8617_out0;
assign v_S_1429_out0 = v_S_9299_out0;
assign v_S_1653_out0 = v_S_9763_out0;
assign v_G1_4205_out0 = v_CARRY_5298_out0 || v_CARRY_5297_out0;
assign v_G1_4429_out0 = v_CARRY_5762_out0 || v_CARRY_5761_out0;
assign v_COUT_897_out0 = v_G1_4205_out0;
assign v_COUT_1121_out0 = v_G1_4429_out0;
assign v__4563_out0 = { v__1839_out0,v_S_1429_out0 };
assign v__4578_out0 = { v__1854_out0,v_S_1653_out0 };
assign v_RM_3566_out0 = v_COUT_897_out0;
assign v_RM_3790_out0 = v_COUT_1121_out0;
assign v_RM_11739_out0 = v_RM_3566_out0;
assign v_RM_12203_out0 = v_RM_3790_out0;
assign v_G1_8154_out0 = ((v_RD_6299_out0 && !v_RM_11739_out0) || (!v_RD_6299_out0) && v_RM_11739_out0);
assign v_G1_8618_out0 = ((v_RD_6763_out0 && !v_RM_12203_out0) || (!v_RD_6763_out0) && v_RM_12203_out0);
assign v_G2_12690_out0 = v_RD_6299_out0 && v_RM_11739_out0;
assign v_G2_13154_out0 = v_RD_6763_out0 && v_RM_12203_out0;
assign v_CARRY_5299_out0 = v_G2_12690_out0;
assign v_CARRY_5763_out0 = v_G2_13154_out0;
assign v_S_9300_out0 = v_G1_8154_out0;
assign v_S_9764_out0 = v_G1_8618_out0;
assign v_RM_11740_out0 = v_S_9300_out0;
assign v_RM_12204_out0 = v_S_9764_out0;
assign v_G1_8155_out0 = ((v_RD_6300_out0 && !v_RM_11740_out0) || (!v_RD_6300_out0) && v_RM_11740_out0);
assign v_G1_8619_out0 = ((v_RD_6764_out0 && !v_RM_12204_out0) || (!v_RD_6764_out0) && v_RM_12204_out0);
assign v_G2_12691_out0 = v_RD_6300_out0 && v_RM_11740_out0;
assign v_G2_13155_out0 = v_RD_6764_out0 && v_RM_12204_out0;
assign v_CARRY_5300_out0 = v_G2_12691_out0;
assign v_CARRY_5764_out0 = v_G2_13155_out0;
assign v_S_9301_out0 = v_G1_8155_out0;
assign v_S_9765_out0 = v_G1_8619_out0;
assign v_S_1430_out0 = v_S_9301_out0;
assign v_S_1654_out0 = v_S_9765_out0;
assign v_G1_4206_out0 = v_CARRY_5300_out0 || v_CARRY_5299_out0;
assign v_G1_4430_out0 = v_CARRY_5764_out0 || v_CARRY_5763_out0;
assign v_COUT_898_out0 = v_G1_4206_out0;
assign v_COUT_1122_out0 = v_G1_4430_out0;
assign v__10665_out0 = { v__4563_out0,v_S_1430_out0 };
assign v__10680_out0 = { v__4578_out0,v_S_1654_out0 };
assign v__10960_out0 = { v__10665_out0,v_COUT_898_out0 };
assign v__10975_out0 = { v__10680_out0,v_COUT_1122_out0 };
assign v_COUT_10930_out0 = v__10960_out0;
assign v_COUT_10945_out0 = v__10975_out0;
assign v_CIN_2360_out0 = v_COUT_10930_out0;
assign v_CIN_2375_out0 = v_COUT_10945_out0;
assign v__473_out0 = v_CIN_2360_out0[8:8];
assign v__488_out0 = v_CIN_2375_out0[8:8];
assign v__1778_out0 = v_CIN_2360_out0[6:6];
assign v__1793_out0 = v_CIN_2375_out0[6:6];
assign v__2160_out0 = v_CIN_2360_out0[3:3];
assign v__2175_out0 = v_CIN_2375_out0[3:3];
assign v__2199_out0 = v_CIN_2360_out0[15:15];
assign v__2213_out0 = v_CIN_2375_out0[15:15];
assign v__2507_out0 = v_CIN_2360_out0[0:0];
assign v__2522_out0 = v_CIN_2375_out0[0:0];
assign v__3056_out0 = v_CIN_2360_out0[9:9];
assign v__3071_out0 = v_CIN_2375_out0[9:9];
assign v__3090_out0 = v_CIN_2360_out0[2:2];
assign v__3105_out0 = v_CIN_2375_out0[2:2];
assign v__3144_out0 = v_CIN_2360_out0[7:7];
assign v__3159_out0 = v_CIN_2375_out0[7:7];
assign v__3828_out0 = v_CIN_2360_out0[1:1];
assign v__3843_out0 = v_CIN_2375_out0[1:1];
assign v__3866_out0 = v_CIN_2360_out0[10:10];
assign v__3881_out0 = v_CIN_2375_out0[10:10];
assign v__6805_out0 = v_CIN_2360_out0[11:11];
assign v__6820_out0 = v_CIN_2375_out0[11:11];
assign v__7649_out0 = v_CIN_2360_out0[12:12];
assign v__7664_out0 = v_CIN_2375_out0[12:12];
assign v__8704_out0 = v_CIN_2360_out0[13:13];
assign v__8719_out0 = v_CIN_2375_out0[13:13];
assign v__8774_out0 = v_CIN_2360_out0[14:14];
assign v__8789_out0 = v_CIN_2375_out0[14:14];
assign v__10724_out0 = v_CIN_2360_out0[5:5];
assign v__10739_out0 = v_CIN_2375_out0[5:5];
assign v__13453_out0 = v_CIN_2360_out0[4:4];
assign v__13468_out0 = v_CIN_2375_out0[4:4];
assign v_RM_3429_out0 = v__7649_out0;
assign v_RM_3430_out0 = v__8774_out0;
assign v_RM_3432_out0 = v__10724_out0;
assign v_RM_3433_out0 = v__13453_out0;
assign v_RM_3434_out0 = v__8704_out0;
assign v_RM_3435_out0 = v__3056_out0;
assign v_RM_3436_out0 = v__3866_out0;
assign v_RM_3437_out0 = v__3828_out0;
assign v_RM_3438_out0 = v__2160_out0;
assign v_RM_3439_out0 = v__1778_out0;
assign v_RM_3440_out0 = v__3144_out0;
assign v_RM_3441_out0 = v__6805_out0;
assign v_RM_3442_out0 = v__473_out0;
assign v_RM_3443_out0 = v__3090_out0;
assign v_RM_3653_out0 = v__7664_out0;
assign v_RM_3654_out0 = v__8789_out0;
assign v_RM_3656_out0 = v__10739_out0;
assign v_RM_3657_out0 = v__13468_out0;
assign v_RM_3658_out0 = v__8719_out0;
assign v_RM_3659_out0 = v__3071_out0;
assign v_RM_3660_out0 = v__3881_out0;
assign v_RM_3661_out0 = v__3843_out0;
assign v_RM_3662_out0 = v__2175_out0;
assign v_RM_3663_out0 = v__1793_out0;
assign v_RM_3664_out0 = v__3159_out0;
assign v_RM_3665_out0 = v__6820_out0;
assign v_RM_3666_out0 = v__488_out0;
assign v_RM_3667_out0 = v__3105_out0;
assign v_CIN_9884_out0 = v__2199_out0;
assign v_CIN_10108_out0 = v__2213_out0;
assign v_RM_11468_out0 = v__2507_out0;
assign v_RM_11932_out0 = v__2522_out0;
assign v_RD_6021_out0 = v_CIN_9884_out0;
assign v_RD_6485_out0 = v_CIN_10108_out0;
assign v_G1_7883_out0 = ((v_RD_6028_out0 && !v_RM_11468_out0) || (!v_RD_6028_out0) && v_RM_11468_out0);
assign v_G1_8347_out0 = ((v_RD_6492_out0 && !v_RM_11932_out0) || (!v_RD_6492_out0) && v_RM_11932_out0);
assign v_RM_11456_out0 = v_RM_3429_out0;
assign v_RM_11458_out0 = v_RM_3430_out0;
assign v_RM_11462_out0 = v_RM_3432_out0;
assign v_RM_11464_out0 = v_RM_3433_out0;
assign v_RM_11466_out0 = v_RM_3434_out0;
assign v_RM_11469_out0 = v_RM_3435_out0;
assign v_RM_11471_out0 = v_RM_3436_out0;
assign v_RM_11473_out0 = v_RM_3437_out0;
assign v_RM_11475_out0 = v_RM_3438_out0;
assign v_RM_11477_out0 = v_RM_3439_out0;
assign v_RM_11479_out0 = v_RM_3440_out0;
assign v_RM_11481_out0 = v_RM_3441_out0;
assign v_RM_11483_out0 = v_RM_3442_out0;
assign v_RM_11485_out0 = v_RM_3443_out0;
assign v_RM_11920_out0 = v_RM_3653_out0;
assign v_RM_11922_out0 = v_RM_3654_out0;
assign v_RM_11926_out0 = v_RM_3656_out0;
assign v_RM_11928_out0 = v_RM_3657_out0;
assign v_RM_11930_out0 = v_RM_3658_out0;
assign v_RM_11933_out0 = v_RM_3659_out0;
assign v_RM_11935_out0 = v_RM_3660_out0;
assign v_RM_11937_out0 = v_RM_3661_out0;
assign v_RM_11939_out0 = v_RM_3662_out0;
assign v_RM_11941_out0 = v_RM_3663_out0;
assign v_RM_11943_out0 = v_RM_3664_out0;
assign v_RM_11945_out0 = v_RM_3665_out0;
assign v_RM_11947_out0 = v_RM_3666_out0;
assign v_RM_11949_out0 = v_RM_3667_out0;
assign v_G2_12419_out0 = v_RD_6028_out0 && v_RM_11468_out0;
assign v_G2_12883_out0 = v_RD_6492_out0 && v_RM_11932_out0;
assign v_CARRY_5028_out0 = v_G2_12419_out0;
assign v_CARRY_5492_out0 = v_G2_12883_out0;
assign v_G1_7871_out0 = ((v_RD_6016_out0 && !v_RM_11456_out0) || (!v_RD_6016_out0) && v_RM_11456_out0);
assign v_G1_7873_out0 = ((v_RD_6018_out0 && !v_RM_11458_out0) || (!v_RD_6018_out0) && v_RM_11458_out0);
assign v_G1_7877_out0 = ((v_RD_6022_out0 && !v_RM_11462_out0) || (!v_RD_6022_out0) && v_RM_11462_out0);
assign v_G1_7879_out0 = ((v_RD_6024_out0 && !v_RM_11464_out0) || (!v_RD_6024_out0) && v_RM_11464_out0);
assign v_G1_7881_out0 = ((v_RD_6026_out0 && !v_RM_11466_out0) || (!v_RD_6026_out0) && v_RM_11466_out0);
assign v_G1_7884_out0 = ((v_RD_6029_out0 && !v_RM_11469_out0) || (!v_RD_6029_out0) && v_RM_11469_out0);
assign v_G1_7886_out0 = ((v_RD_6031_out0 && !v_RM_11471_out0) || (!v_RD_6031_out0) && v_RM_11471_out0);
assign v_G1_7888_out0 = ((v_RD_6033_out0 && !v_RM_11473_out0) || (!v_RD_6033_out0) && v_RM_11473_out0);
assign v_G1_7890_out0 = ((v_RD_6035_out0 && !v_RM_11475_out0) || (!v_RD_6035_out0) && v_RM_11475_out0);
assign v_G1_7892_out0 = ((v_RD_6037_out0 && !v_RM_11477_out0) || (!v_RD_6037_out0) && v_RM_11477_out0);
assign v_G1_7894_out0 = ((v_RD_6039_out0 && !v_RM_11479_out0) || (!v_RD_6039_out0) && v_RM_11479_out0);
assign v_G1_7896_out0 = ((v_RD_6041_out0 && !v_RM_11481_out0) || (!v_RD_6041_out0) && v_RM_11481_out0);
assign v_G1_7898_out0 = ((v_RD_6043_out0 && !v_RM_11483_out0) || (!v_RD_6043_out0) && v_RM_11483_out0);
assign v_G1_7900_out0 = ((v_RD_6045_out0 && !v_RM_11485_out0) || (!v_RD_6045_out0) && v_RM_11485_out0);
assign v_G1_8335_out0 = ((v_RD_6480_out0 && !v_RM_11920_out0) || (!v_RD_6480_out0) && v_RM_11920_out0);
assign v_G1_8337_out0 = ((v_RD_6482_out0 && !v_RM_11922_out0) || (!v_RD_6482_out0) && v_RM_11922_out0);
assign v_G1_8341_out0 = ((v_RD_6486_out0 && !v_RM_11926_out0) || (!v_RD_6486_out0) && v_RM_11926_out0);
assign v_G1_8343_out0 = ((v_RD_6488_out0 && !v_RM_11928_out0) || (!v_RD_6488_out0) && v_RM_11928_out0);
assign v_G1_8345_out0 = ((v_RD_6490_out0 && !v_RM_11930_out0) || (!v_RD_6490_out0) && v_RM_11930_out0);
assign v_G1_8348_out0 = ((v_RD_6493_out0 && !v_RM_11933_out0) || (!v_RD_6493_out0) && v_RM_11933_out0);
assign v_G1_8350_out0 = ((v_RD_6495_out0 && !v_RM_11935_out0) || (!v_RD_6495_out0) && v_RM_11935_out0);
assign v_G1_8352_out0 = ((v_RD_6497_out0 && !v_RM_11937_out0) || (!v_RD_6497_out0) && v_RM_11937_out0);
assign v_G1_8354_out0 = ((v_RD_6499_out0 && !v_RM_11939_out0) || (!v_RD_6499_out0) && v_RM_11939_out0);
assign v_G1_8356_out0 = ((v_RD_6501_out0 && !v_RM_11941_out0) || (!v_RD_6501_out0) && v_RM_11941_out0);
assign v_G1_8358_out0 = ((v_RD_6503_out0 && !v_RM_11943_out0) || (!v_RD_6503_out0) && v_RM_11943_out0);
assign v_G1_8360_out0 = ((v_RD_6505_out0 && !v_RM_11945_out0) || (!v_RD_6505_out0) && v_RM_11945_out0);
assign v_G1_8362_out0 = ((v_RD_6507_out0 && !v_RM_11947_out0) || (!v_RD_6507_out0) && v_RM_11947_out0);
assign v_G1_8364_out0 = ((v_RD_6509_out0 && !v_RM_11949_out0) || (!v_RD_6509_out0) && v_RM_11949_out0);
assign v_S_9029_out0 = v_G1_7883_out0;
assign v_S_9493_out0 = v_G1_8347_out0;
assign v_G2_12407_out0 = v_RD_6016_out0 && v_RM_11456_out0;
assign v_G2_12409_out0 = v_RD_6018_out0 && v_RM_11458_out0;
assign v_G2_12413_out0 = v_RD_6022_out0 && v_RM_11462_out0;
assign v_G2_12415_out0 = v_RD_6024_out0 && v_RM_11464_out0;
assign v_G2_12417_out0 = v_RD_6026_out0 && v_RM_11466_out0;
assign v_G2_12420_out0 = v_RD_6029_out0 && v_RM_11469_out0;
assign v_G2_12422_out0 = v_RD_6031_out0 && v_RM_11471_out0;
assign v_G2_12424_out0 = v_RD_6033_out0 && v_RM_11473_out0;
assign v_G2_12426_out0 = v_RD_6035_out0 && v_RM_11475_out0;
assign v_G2_12428_out0 = v_RD_6037_out0 && v_RM_11477_out0;
assign v_G2_12430_out0 = v_RD_6039_out0 && v_RM_11479_out0;
assign v_G2_12432_out0 = v_RD_6041_out0 && v_RM_11481_out0;
assign v_G2_12434_out0 = v_RD_6043_out0 && v_RM_11483_out0;
assign v_G2_12436_out0 = v_RD_6045_out0 && v_RM_11485_out0;
assign v_G2_12871_out0 = v_RD_6480_out0 && v_RM_11920_out0;
assign v_G2_12873_out0 = v_RD_6482_out0 && v_RM_11922_out0;
assign v_G2_12877_out0 = v_RD_6486_out0 && v_RM_11926_out0;
assign v_G2_12879_out0 = v_RD_6488_out0 && v_RM_11928_out0;
assign v_G2_12881_out0 = v_RD_6490_out0 && v_RM_11930_out0;
assign v_G2_12884_out0 = v_RD_6493_out0 && v_RM_11933_out0;
assign v_G2_12886_out0 = v_RD_6495_out0 && v_RM_11935_out0;
assign v_G2_12888_out0 = v_RD_6497_out0 && v_RM_11937_out0;
assign v_G2_12890_out0 = v_RD_6499_out0 && v_RM_11939_out0;
assign v_G2_12892_out0 = v_RD_6501_out0 && v_RM_11941_out0;
assign v_G2_12894_out0 = v_RD_6503_out0 && v_RM_11943_out0;
assign v_G2_12896_out0 = v_RD_6505_out0 && v_RM_11945_out0;
assign v_G2_12898_out0 = v_RD_6507_out0 && v_RM_11947_out0;
assign v_G2_12900_out0 = v_RD_6509_out0 && v_RM_11949_out0;
assign v_S_4670_out0 = v_S_9029_out0;
assign v_S_4685_out0 = v_S_9493_out0;
assign v_CARRY_5016_out0 = v_G2_12407_out0;
assign v_CARRY_5018_out0 = v_G2_12409_out0;
assign v_CARRY_5022_out0 = v_G2_12413_out0;
assign v_CARRY_5024_out0 = v_G2_12415_out0;
assign v_CARRY_5026_out0 = v_G2_12417_out0;
assign v_CARRY_5029_out0 = v_G2_12420_out0;
assign v_CARRY_5031_out0 = v_G2_12422_out0;
assign v_CARRY_5033_out0 = v_G2_12424_out0;
assign v_CARRY_5035_out0 = v_G2_12426_out0;
assign v_CARRY_5037_out0 = v_G2_12428_out0;
assign v_CARRY_5039_out0 = v_G2_12430_out0;
assign v_CARRY_5041_out0 = v_G2_12432_out0;
assign v_CARRY_5043_out0 = v_G2_12434_out0;
assign v_CARRY_5045_out0 = v_G2_12436_out0;
assign v_CARRY_5480_out0 = v_G2_12871_out0;
assign v_CARRY_5482_out0 = v_G2_12873_out0;
assign v_CARRY_5486_out0 = v_G2_12877_out0;
assign v_CARRY_5488_out0 = v_G2_12879_out0;
assign v_CARRY_5490_out0 = v_G2_12881_out0;
assign v_CARRY_5493_out0 = v_G2_12884_out0;
assign v_CARRY_5495_out0 = v_G2_12886_out0;
assign v_CARRY_5497_out0 = v_G2_12888_out0;
assign v_CARRY_5499_out0 = v_G2_12890_out0;
assign v_CARRY_5501_out0 = v_G2_12892_out0;
assign v_CARRY_5503_out0 = v_G2_12894_out0;
assign v_CARRY_5505_out0 = v_G2_12896_out0;
assign v_CARRY_5507_out0 = v_G2_12898_out0;
assign v_CARRY_5509_out0 = v_G2_12900_out0;
assign v_S_9017_out0 = v_G1_7871_out0;
assign v_S_9019_out0 = v_G1_7873_out0;
assign v_S_9023_out0 = v_G1_7877_out0;
assign v_S_9025_out0 = v_G1_7879_out0;
assign v_S_9027_out0 = v_G1_7881_out0;
assign v_S_9030_out0 = v_G1_7884_out0;
assign v_S_9032_out0 = v_G1_7886_out0;
assign v_S_9034_out0 = v_G1_7888_out0;
assign v_S_9036_out0 = v_G1_7890_out0;
assign v_S_9038_out0 = v_G1_7892_out0;
assign v_S_9040_out0 = v_G1_7894_out0;
assign v_S_9042_out0 = v_G1_7896_out0;
assign v_S_9044_out0 = v_G1_7898_out0;
assign v_S_9046_out0 = v_G1_7900_out0;
assign v_S_9481_out0 = v_G1_8335_out0;
assign v_S_9483_out0 = v_G1_8337_out0;
assign v_S_9487_out0 = v_G1_8341_out0;
assign v_S_9489_out0 = v_G1_8343_out0;
assign v_S_9491_out0 = v_G1_8345_out0;
assign v_S_9494_out0 = v_G1_8348_out0;
assign v_S_9496_out0 = v_G1_8350_out0;
assign v_S_9498_out0 = v_G1_8352_out0;
assign v_S_9500_out0 = v_G1_8354_out0;
assign v_S_9502_out0 = v_G1_8356_out0;
assign v_S_9504_out0 = v_G1_8358_out0;
assign v_S_9506_out0 = v_G1_8360_out0;
assign v_S_9508_out0 = v_G1_8362_out0;
assign v_S_9510_out0 = v_G1_8364_out0;
assign v_CIN_9890_out0 = v_CARRY_5028_out0;
assign v_CIN_10114_out0 = v_CARRY_5492_out0;
assign v__2191_out0 = { v__10775_out0,v_S_4670_out0 };
assign v__2192_out0 = { v__10776_out0,v_S_4685_out0 };
assign v_RD_6034_out0 = v_CIN_9890_out0;
assign v_RD_6498_out0 = v_CIN_10114_out0;
assign v_RM_11457_out0 = v_S_9017_out0;
assign v_RM_11459_out0 = v_S_9019_out0;
assign v_RM_11463_out0 = v_S_9023_out0;
assign v_RM_11465_out0 = v_S_9025_out0;
assign v_RM_11467_out0 = v_S_9027_out0;
assign v_RM_11470_out0 = v_S_9030_out0;
assign v_RM_11472_out0 = v_S_9032_out0;
assign v_RM_11474_out0 = v_S_9034_out0;
assign v_RM_11476_out0 = v_S_9036_out0;
assign v_RM_11478_out0 = v_S_9038_out0;
assign v_RM_11480_out0 = v_S_9040_out0;
assign v_RM_11482_out0 = v_S_9042_out0;
assign v_RM_11484_out0 = v_S_9044_out0;
assign v_RM_11486_out0 = v_S_9046_out0;
assign v_RM_11921_out0 = v_S_9481_out0;
assign v_RM_11923_out0 = v_S_9483_out0;
assign v_RM_11927_out0 = v_S_9487_out0;
assign v_RM_11929_out0 = v_S_9489_out0;
assign v_RM_11931_out0 = v_S_9491_out0;
assign v_RM_11934_out0 = v_S_9494_out0;
assign v_RM_11936_out0 = v_S_9496_out0;
assign v_RM_11938_out0 = v_S_9498_out0;
assign v_RM_11940_out0 = v_S_9500_out0;
assign v_RM_11942_out0 = v_S_9502_out0;
assign v_RM_11944_out0 = v_S_9504_out0;
assign v_RM_11946_out0 = v_S_9506_out0;
assign v_RM_11948_out0 = v_S_9508_out0;
assign v_RM_11950_out0 = v_S_9510_out0;
assign v_G1_7889_out0 = ((v_RD_6034_out0 && !v_RM_11474_out0) || (!v_RD_6034_out0) && v_RM_11474_out0);
assign v_G1_8353_out0 = ((v_RD_6498_out0 && !v_RM_11938_out0) || (!v_RD_6498_out0) && v_RM_11938_out0);
assign v_G2_12425_out0 = v_RD_6034_out0 && v_RM_11474_out0;
assign v_G2_12889_out0 = v_RD_6498_out0 && v_RM_11938_out0;
assign v_CARRY_5034_out0 = v_G2_12425_out0;
assign v_CARRY_5498_out0 = v_G2_12889_out0;
assign v_S_9035_out0 = v_G1_7889_out0;
assign v_S_9499_out0 = v_G1_8353_out0;
assign v_S_1301_out0 = v_S_9035_out0;
assign v_S_1525_out0 = v_S_9499_out0;
assign v_G1_4077_out0 = v_CARRY_5034_out0 || v_CARRY_5033_out0;
assign v_G1_4301_out0 = v_CARRY_5498_out0 || v_CARRY_5497_out0;
assign v_COUT_769_out0 = v_G1_4077_out0;
assign v_COUT_993_out0 = v_G1_4301_out0;
assign v_CIN_9896_out0 = v_COUT_769_out0;
assign v_CIN_10120_out0 = v_COUT_993_out0;
assign v_RD_6046_out0 = v_CIN_9896_out0;
assign v_RD_6510_out0 = v_CIN_10120_out0;
assign v_G1_7901_out0 = ((v_RD_6046_out0 && !v_RM_11486_out0) || (!v_RD_6046_out0) && v_RM_11486_out0);
assign v_G1_8365_out0 = ((v_RD_6510_out0 && !v_RM_11950_out0) || (!v_RD_6510_out0) && v_RM_11950_out0);
assign v_G2_12437_out0 = v_RD_6046_out0 && v_RM_11486_out0;
assign v_G2_12901_out0 = v_RD_6510_out0 && v_RM_11950_out0;
assign v_CARRY_5046_out0 = v_G2_12437_out0;
assign v_CARRY_5510_out0 = v_G2_12901_out0;
assign v_S_9047_out0 = v_G1_7901_out0;
assign v_S_9511_out0 = v_G1_8365_out0;
assign v_S_1307_out0 = v_S_9047_out0;
assign v_S_1531_out0 = v_S_9511_out0;
assign v_G1_4083_out0 = v_CARRY_5046_out0 || v_CARRY_5045_out0;
assign v_G1_4307_out0 = v_CARRY_5510_out0 || v_CARRY_5509_out0;
assign v_COUT_775_out0 = v_G1_4083_out0;
assign v_COUT_999_out0 = v_G1_4307_out0;
assign v__4787_out0 = { v_S_1301_out0,v_S_1307_out0 };
assign v__4802_out0 = { v_S_1525_out0,v_S_1531_out0 };
assign v_CIN_9891_out0 = v_COUT_775_out0;
assign v_CIN_10115_out0 = v_COUT_999_out0;
assign v_RD_6036_out0 = v_CIN_9891_out0;
assign v_RD_6500_out0 = v_CIN_10115_out0;
assign v_G1_7891_out0 = ((v_RD_6036_out0 && !v_RM_11476_out0) || (!v_RD_6036_out0) && v_RM_11476_out0);
assign v_G1_8355_out0 = ((v_RD_6500_out0 && !v_RM_11940_out0) || (!v_RD_6500_out0) && v_RM_11940_out0);
assign v_G2_12427_out0 = v_RD_6036_out0 && v_RM_11476_out0;
assign v_G2_12891_out0 = v_RD_6500_out0 && v_RM_11940_out0;
assign v_CARRY_5036_out0 = v_G2_12427_out0;
assign v_CARRY_5500_out0 = v_G2_12891_out0;
assign v_S_9037_out0 = v_G1_7891_out0;
assign v_S_9501_out0 = v_G1_8355_out0;
assign v_S_1302_out0 = v_S_9037_out0;
assign v_S_1526_out0 = v_S_9501_out0;
assign v_G1_4078_out0 = v_CARRY_5036_out0 || v_CARRY_5035_out0;
assign v_G1_4302_out0 = v_CARRY_5500_out0 || v_CARRY_5499_out0;
assign v_COUT_770_out0 = v_G1_4078_out0;
assign v_COUT_994_out0 = v_G1_4302_out0;
assign v__2557_out0 = { v__4787_out0,v_S_1302_out0 };
assign v__2572_out0 = { v__4802_out0,v_S_1526_out0 };
assign v_CIN_9886_out0 = v_COUT_770_out0;
assign v_CIN_10110_out0 = v_COUT_994_out0;
assign v_RD_6025_out0 = v_CIN_9886_out0;
assign v_RD_6489_out0 = v_CIN_10110_out0;
assign v_G1_7880_out0 = ((v_RD_6025_out0 && !v_RM_11465_out0) || (!v_RD_6025_out0) && v_RM_11465_out0);
assign v_G1_8344_out0 = ((v_RD_6489_out0 && !v_RM_11929_out0) || (!v_RD_6489_out0) && v_RM_11929_out0);
assign v_G2_12416_out0 = v_RD_6025_out0 && v_RM_11465_out0;
assign v_G2_12880_out0 = v_RD_6489_out0 && v_RM_11929_out0;
assign v_CARRY_5025_out0 = v_G2_12416_out0;
assign v_CARRY_5489_out0 = v_G2_12880_out0;
assign v_S_9026_out0 = v_G1_7880_out0;
assign v_S_9490_out0 = v_G1_8344_out0;
assign v_S_1297_out0 = v_S_9026_out0;
assign v_S_1521_out0 = v_S_9490_out0;
assign v_G1_4073_out0 = v_CARRY_5025_out0 || v_CARRY_5024_out0;
assign v_G1_4297_out0 = v_CARRY_5489_out0 || v_CARRY_5488_out0;
assign v_COUT_765_out0 = v_G1_4073_out0;
assign v_COUT_989_out0 = v_G1_4297_out0;
assign v__7037_out0 = { v__2557_out0,v_S_1297_out0 };
assign v__7052_out0 = { v__2572_out0,v_S_1521_out0 };
assign v_CIN_9885_out0 = v_COUT_765_out0;
assign v_CIN_10109_out0 = v_COUT_989_out0;
assign v_RD_6023_out0 = v_CIN_9885_out0;
assign v_RD_6487_out0 = v_CIN_10109_out0;
assign v_G1_7878_out0 = ((v_RD_6023_out0 && !v_RM_11463_out0) || (!v_RD_6023_out0) && v_RM_11463_out0);
assign v_G1_8342_out0 = ((v_RD_6487_out0 && !v_RM_11927_out0) || (!v_RD_6487_out0) && v_RM_11927_out0);
assign v_G2_12414_out0 = v_RD_6023_out0 && v_RM_11463_out0;
assign v_G2_12878_out0 = v_RD_6487_out0 && v_RM_11927_out0;
assign v_CARRY_5023_out0 = v_G2_12414_out0;
assign v_CARRY_5487_out0 = v_G2_12878_out0;
assign v_S_9024_out0 = v_G1_7878_out0;
assign v_S_9488_out0 = v_G1_8342_out0;
assign v_S_1296_out0 = v_S_9024_out0;
assign v_S_1520_out0 = v_S_9488_out0;
assign v_G1_4072_out0 = v_CARRY_5023_out0 || v_CARRY_5022_out0;
assign v_G1_4296_out0 = v_CARRY_5487_out0 || v_CARRY_5486_out0;
assign v_COUT_764_out0 = v_G1_4072_out0;
assign v_COUT_988_out0 = v_G1_4296_out0;
assign v__13523_out0 = { v__7037_out0,v_S_1296_out0 };
assign v__13538_out0 = { v__7052_out0,v_S_1520_out0 };
assign v_CIN_9892_out0 = v_COUT_764_out0;
assign v_CIN_10116_out0 = v_COUT_988_out0;
assign v_RD_6038_out0 = v_CIN_9892_out0;
assign v_RD_6502_out0 = v_CIN_10116_out0;
assign v_G1_7893_out0 = ((v_RD_6038_out0 && !v_RM_11478_out0) || (!v_RD_6038_out0) && v_RM_11478_out0);
assign v_G1_8357_out0 = ((v_RD_6502_out0 && !v_RM_11942_out0) || (!v_RD_6502_out0) && v_RM_11942_out0);
assign v_G2_12429_out0 = v_RD_6038_out0 && v_RM_11478_out0;
assign v_G2_12893_out0 = v_RD_6502_out0 && v_RM_11942_out0;
assign v_CARRY_5038_out0 = v_G2_12429_out0;
assign v_CARRY_5502_out0 = v_G2_12893_out0;
assign v_S_9039_out0 = v_G1_7893_out0;
assign v_S_9503_out0 = v_G1_8357_out0;
assign v_S_1303_out0 = v_S_9039_out0;
assign v_S_1527_out0 = v_S_9503_out0;
assign v_G1_4079_out0 = v_CARRY_5038_out0 || v_CARRY_5037_out0;
assign v_G1_4303_out0 = v_CARRY_5502_out0 || v_CARRY_5501_out0;
assign v_COUT_771_out0 = v_G1_4079_out0;
assign v_COUT_995_out0 = v_G1_4303_out0;
assign v__3316_out0 = { v__13523_out0,v_S_1303_out0 };
assign v__3331_out0 = { v__13538_out0,v_S_1527_out0 };
assign v_CIN_9893_out0 = v_COUT_771_out0;
assign v_CIN_10117_out0 = v_COUT_995_out0;
assign v_RD_6040_out0 = v_CIN_9893_out0;
assign v_RD_6504_out0 = v_CIN_10117_out0;
assign v_G1_7895_out0 = ((v_RD_6040_out0 && !v_RM_11480_out0) || (!v_RD_6040_out0) && v_RM_11480_out0);
assign v_G1_8359_out0 = ((v_RD_6504_out0 && !v_RM_11944_out0) || (!v_RD_6504_out0) && v_RM_11944_out0);
assign v_G2_12431_out0 = v_RD_6040_out0 && v_RM_11480_out0;
assign v_G2_12895_out0 = v_RD_6504_out0 && v_RM_11944_out0;
assign v_CARRY_5040_out0 = v_G2_12431_out0;
assign v_CARRY_5504_out0 = v_G2_12895_out0;
assign v_S_9041_out0 = v_G1_7895_out0;
assign v_S_9505_out0 = v_G1_8359_out0;
assign v_S_1304_out0 = v_S_9041_out0;
assign v_S_1528_out0 = v_S_9505_out0;
assign v_G1_4080_out0 = v_CARRY_5040_out0 || v_CARRY_5039_out0;
assign v_G1_4304_out0 = v_CARRY_5504_out0 || v_CARRY_5503_out0;
assign v_COUT_772_out0 = v_G1_4080_out0;
assign v_COUT_996_out0 = v_G1_4304_out0;
assign v__7152_out0 = { v__3316_out0,v_S_1304_out0 };
assign v__7167_out0 = { v__3331_out0,v_S_1528_out0 };
assign v_CIN_9895_out0 = v_COUT_772_out0;
assign v_CIN_10119_out0 = v_COUT_996_out0;
assign v_RD_6044_out0 = v_CIN_9895_out0;
assign v_RD_6508_out0 = v_CIN_10119_out0;
assign v_G1_7899_out0 = ((v_RD_6044_out0 && !v_RM_11484_out0) || (!v_RD_6044_out0) && v_RM_11484_out0);
assign v_G1_8363_out0 = ((v_RD_6508_out0 && !v_RM_11948_out0) || (!v_RD_6508_out0) && v_RM_11948_out0);
assign v_G2_12435_out0 = v_RD_6044_out0 && v_RM_11484_out0;
assign v_G2_12899_out0 = v_RD_6508_out0 && v_RM_11948_out0;
assign v_CARRY_5044_out0 = v_G2_12435_out0;
assign v_CARRY_5508_out0 = v_G2_12899_out0;
assign v_S_9045_out0 = v_G1_7899_out0;
assign v_S_9509_out0 = v_G1_8363_out0;
assign v_S_1306_out0 = v_S_9045_out0;
assign v_S_1530_out0 = v_S_9509_out0;
assign v_G1_4082_out0 = v_CARRY_5044_out0 || v_CARRY_5043_out0;
assign v_G1_4306_out0 = v_CARRY_5508_out0 || v_CARRY_5507_out0;
assign v_COUT_774_out0 = v_G1_4082_out0;
assign v_COUT_998_out0 = v_G1_4306_out0;
assign v__4754_out0 = { v__7152_out0,v_S_1306_out0 };
assign v__4769_out0 = { v__7167_out0,v_S_1530_out0 };
assign v_CIN_9888_out0 = v_COUT_774_out0;
assign v_CIN_10112_out0 = v_COUT_998_out0;
assign v_RD_6030_out0 = v_CIN_9888_out0;
assign v_RD_6494_out0 = v_CIN_10112_out0;
assign v_G1_7885_out0 = ((v_RD_6030_out0 && !v_RM_11470_out0) || (!v_RD_6030_out0) && v_RM_11470_out0);
assign v_G1_8349_out0 = ((v_RD_6494_out0 && !v_RM_11934_out0) || (!v_RD_6494_out0) && v_RM_11934_out0);
assign v_G2_12421_out0 = v_RD_6030_out0 && v_RM_11470_out0;
assign v_G2_12885_out0 = v_RD_6494_out0 && v_RM_11934_out0;
assign v_CARRY_5030_out0 = v_G2_12421_out0;
assign v_CARRY_5494_out0 = v_G2_12885_out0;
assign v_S_9031_out0 = v_G1_7885_out0;
assign v_S_9495_out0 = v_G1_8349_out0;
assign v_S_1299_out0 = v_S_9031_out0;
assign v_S_1523_out0 = v_S_9495_out0;
assign v_G1_4075_out0 = v_CARRY_5030_out0 || v_CARRY_5029_out0;
assign v_G1_4299_out0 = v_CARRY_5494_out0 || v_CARRY_5493_out0;
assign v_COUT_767_out0 = v_G1_4075_out0;
assign v_COUT_991_out0 = v_G1_4299_out0;
assign v__6931_out0 = { v__4754_out0,v_S_1299_out0 };
assign v__6946_out0 = { v__4769_out0,v_S_1523_out0 };
assign v_CIN_9889_out0 = v_COUT_767_out0;
assign v_CIN_10113_out0 = v_COUT_991_out0;
assign v_RD_6032_out0 = v_CIN_9889_out0;
assign v_RD_6496_out0 = v_CIN_10113_out0;
assign v_G1_7887_out0 = ((v_RD_6032_out0 && !v_RM_11472_out0) || (!v_RD_6032_out0) && v_RM_11472_out0);
assign v_G1_8351_out0 = ((v_RD_6496_out0 && !v_RM_11936_out0) || (!v_RD_6496_out0) && v_RM_11936_out0);
assign v_G2_12423_out0 = v_RD_6032_out0 && v_RM_11472_out0;
assign v_G2_12887_out0 = v_RD_6496_out0 && v_RM_11936_out0;
assign v_CARRY_5032_out0 = v_G2_12423_out0;
assign v_CARRY_5496_out0 = v_G2_12887_out0;
assign v_S_9033_out0 = v_G1_7887_out0;
assign v_S_9497_out0 = v_G1_8351_out0;
assign v_S_1300_out0 = v_S_9033_out0;
assign v_S_1524_out0 = v_S_9497_out0;
assign v_G1_4076_out0 = v_CARRY_5032_out0 || v_CARRY_5031_out0;
assign v_G1_4300_out0 = v_CARRY_5496_out0 || v_CARRY_5495_out0;
assign v_COUT_768_out0 = v_G1_4076_out0;
assign v_COUT_992_out0 = v_G1_4300_out0;
assign v__5807_out0 = { v__6931_out0,v_S_1300_out0 };
assign v__5822_out0 = { v__6946_out0,v_S_1524_out0 };
assign v_CIN_9894_out0 = v_COUT_768_out0;
assign v_CIN_10118_out0 = v_COUT_992_out0;
assign v_RD_6042_out0 = v_CIN_9894_out0;
assign v_RD_6506_out0 = v_CIN_10118_out0;
assign v_G1_7897_out0 = ((v_RD_6042_out0 && !v_RM_11482_out0) || (!v_RD_6042_out0) && v_RM_11482_out0);
assign v_G1_8361_out0 = ((v_RD_6506_out0 && !v_RM_11946_out0) || (!v_RD_6506_out0) && v_RM_11946_out0);
assign v_G2_12433_out0 = v_RD_6042_out0 && v_RM_11482_out0;
assign v_G2_12897_out0 = v_RD_6506_out0 && v_RM_11946_out0;
assign v_CARRY_5042_out0 = v_G2_12433_out0;
assign v_CARRY_5506_out0 = v_G2_12897_out0;
assign v_S_9043_out0 = v_G1_7897_out0;
assign v_S_9507_out0 = v_G1_8361_out0;
assign v_S_1305_out0 = v_S_9043_out0;
assign v_S_1529_out0 = v_S_9507_out0;
assign v_G1_4081_out0 = v_CARRY_5042_out0 || v_CARRY_5041_out0;
assign v_G1_4305_out0 = v_CARRY_5506_out0 || v_CARRY_5505_out0;
assign v_COUT_773_out0 = v_G1_4081_out0;
assign v_COUT_997_out0 = v_G1_4305_out0;
assign v__2031_out0 = { v__5807_out0,v_S_1305_out0 };
assign v__2046_out0 = { v__5822_out0,v_S_1529_out0 };
assign v_CIN_9882_out0 = v_COUT_773_out0;
assign v_CIN_10106_out0 = v_COUT_997_out0;
assign v_RD_6017_out0 = v_CIN_9882_out0;
assign v_RD_6481_out0 = v_CIN_10106_out0;
assign v_G1_7872_out0 = ((v_RD_6017_out0 && !v_RM_11457_out0) || (!v_RD_6017_out0) && v_RM_11457_out0);
assign v_G1_8336_out0 = ((v_RD_6481_out0 && !v_RM_11921_out0) || (!v_RD_6481_out0) && v_RM_11921_out0);
assign v_G2_12408_out0 = v_RD_6017_out0 && v_RM_11457_out0;
assign v_G2_12872_out0 = v_RD_6481_out0 && v_RM_11921_out0;
assign v_CARRY_5017_out0 = v_G2_12408_out0;
assign v_CARRY_5481_out0 = v_G2_12872_out0;
assign v_S_9018_out0 = v_G1_7872_out0;
assign v_S_9482_out0 = v_G1_8336_out0;
assign v_S_1293_out0 = v_S_9018_out0;
assign v_S_1517_out0 = v_S_9482_out0;
assign v_G1_4069_out0 = v_CARRY_5017_out0 || v_CARRY_5016_out0;
assign v_G1_4293_out0 = v_CARRY_5481_out0 || v_CARRY_5480_out0;
assign v_COUT_761_out0 = v_G1_4069_out0;
assign v_COUT_985_out0 = v_G1_4293_out0;
assign v__2798_out0 = { v__2031_out0,v_S_1293_out0 };
assign v__2813_out0 = { v__2046_out0,v_S_1517_out0 };
assign v_CIN_9887_out0 = v_COUT_761_out0;
assign v_CIN_10111_out0 = v_COUT_985_out0;
assign v_RD_6027_out0 = v_CIN_9887_out0;
assign v_RD_6491_out0 = v_CIN_10111_out0;
assign v_G1_7882_out0 = ((v_RD_6027_out0 && !v_RM_11467_out0) || (!v_RD_6027_out0) && v_RM_11467_out0);
assign v_G1_8346_out0 = ((v_RD_6491_out0 && !v_RM_11931_out0) || (!v_RD_6491_out0) && v_RM_11931_out0);
assign v_G2_12418_out0 = v_RD_6027_out0 && v_RM_11467_out0;
assign v_G2_12882_out0 = v_RD_6491_out0 && v_RM_11931_out0;
assign v_CARRY_5027_out0 = v_G2_12418_out0;
assign v_CARRY_5491_out0 = v_G2_12882_out0;
assign v_S_9028_out0 = v_G1_7882_out0;
assign v_S_9492_out0 = v_G1_8346_out0;
assign v_S_1298_out0 = v_S_9028_out0;
assign v_S_1522_out0 = v_S_9492_out0;
assign v_G1_4074_out0 = v_CARRY_5027_out0 || v_CARRY_5026_out0;
assign v_G1_4298_out0 = v_CARRY_5491_out0 || v_CARRY_5490_out0;
assign v_COUT_766_out0 = v_G1_4074_out0;
assign v_COUT_990_out0 = v_G1_4298_out0;
assign v__1830_out0 = { v__2798_out0,v_S_1298_out0 };
assign v__1845_out0 = { v__2813_out0,v_S_1522_out0 };
assign v_CIN_9883_out0 = v_COUT_766_out0;
assign v_CIN_10107_out0 = v_COUT_990_out0;
assign v_RD_6019_out0 = v_CIN_9883_out0;
assign v_RD_6483_out0 = v_CIN_10107_out0;
assign v_G1_7874_out0 = ((v_RD_6019_out0 && !v_RM_11459_out0) || (!v_RD_6019_out0) && v_RM_11459_out0);
assign v_G1_8338_out0 = ((v_RD_6483_out0 && !v_RM_11923_out0) || (!v_RD_6483_out0) && v_RM_11923_out0);
assign v_G2_12410_out0 = v_RD_6019_out0 && v_RM_11459_out0;
assign v_G2_12874_out0 = v_RD_6483_out0 && v_RM_11923_out0;
assign v_CARRY_5019_out0 = v_G2_12410_out0;
assign v_CARRY_5483_out0 = v_G2_12874_out0;
assign v_S_9020_out0 = v_G1_7874_out0;
assign v_S_9484_out0 = v_G1_8338_out0;
assign v_S_1294_out0 = v_S_9020_out0;
assign v_S_1518_out0 = v_S_9484_out0;
assign v_G1_4070_out0 = v_CARRY_5019_out0 || v_CARRY_5018_out0;
assign v_G1_4294_out0 = v_CARRY_5483_out0 || v_CARRY_5482_out0;
assign v_COUT_762_out0 = v_G1_4070_out0;
assign v_COUT_986_out0 = v_G1_4294_out0;
assign v__4554_out0 = { v__1830_out0,v_S_1294_out0 };
assign v__4569_out0 = { v__1845_out0,v_S_1518_out0 };
assign v_RM_3431_out0 = v_COUT_762_out0;
assign v_RM_3655_out0 = v_COUT_986_out0;
assign v_RM_11460_out0 = v_RM_3431_out0;
assign v_RM_11924_out0 = v_RM_3655_out0;
assign v_G1_7875_out0 = ((v_RD_6020_out0 && !v_RM_11460_out0) || (!v_RD_6020_out0) && v_RM_11460_out0);
assign v_G1_8339_out0 = ((v_RD_6484_out0 && !v_RM_11924_out0) || (!v_RD_6484_out0) && v_RM_11924_out0);
assign v_G2_12411_out0 = v_RD_6020_out0 && v_RM_11460_out0;
assign v_G2_12875_out0 = v_RD_6484_out0 && v_RM_11924_out0;
assign v_CARRY_5020_out0 = v_G2_12411_out0;
assign v_CARRY_5484_out0 = v_G2_12875_out0;
assign v_S_9021_out0 = v_G1_7875_out0;
assign v_S_9485_out0 = v_G1_8339_out0;
assign v_RM_11461_out0 = v_S_9021_out0;
assign v_RM_11925_out0 = v_S_9485_out0;
assign v_G1_7876_out0 = ((v_RD_6021_out0 && !v_RM_11461_out0) || (!v_RD_6021_out0) && v_RM_11461_out0);
assign v_G1_8340_out0 = ((v_RD_6485_out0 && !v_RM_11925_out0) || (!v_RD_6485_out0) && v_RM_11925_out0);
assign v_G2_12412_out0 = v_RD_6021_out0 && v_RM_11461_out0;
assign v_G2_12876_out0 = v_RD_6485_out0 && v_RM_11925_out0;
assign v_CARRY_5021_out0 = v_G2_12412_out0;
assign v_CARRY_5485_out0 = v_G2_12876_out0;
assign v_S_9022_out0 = v_G1_7876_out0;
assign v_S_9486_out0 = v_G1_8340_out0;
assign v_S_1295_out0 = v_S_9022_out0;
assign v_S_1519_out0 = v_S_9486_out0;
assign v_G1_4071_out0 = v_CARRY_5021_out0 || v_CARRY_5020_out0;
assign v_G1_4295_out0 = v_CARRY_5485_out0 || v_CARRY_5484_out0;
assign v_COUT_763_out0 = v_G1_4071_out0;
assign v_COUT_987_out0 = v_G1_4295_out0;
assign v__10656_out0 = { v__4554_out0,v_S_1295_out0 };
assign v__10671_out0 = { v__4569_out0,v_S_1519_out0 };
assign v__10951_out0 = { v__10656_out0,v_COUT_763_out0 };
assign v__10966_out0 = { v__10671_out0,v_COUT_987_out0 };
assign v_COUT_10921_out0 = v__10951_out0;
assign v_COUT_10936_out0 = v__10966_out0;
assign v_CIN_2358_out0 = v_COUT_10921_out0;
assign v_CIN_2373_out0 = v_COUT_10936_out0;
assign v__471_out0 = v_CIN_2358_out0[8:8];
assign v__486_out0 = v_CIN_2373_out0[8:8];
assign v__1776_out0 = v_CIN_2358_out0[6:6];
assign v__1791_out0 = v_CIN_2373_out0[6:6];
assign v__2158_out0 = v_CIN_2358_out0[3:3];
assign v__2173_out0 = v_CIN_2373_out0[3:3];
assign v__2197_out0 = v_CIN_2358_out0[15:15];
assign v__2211_out0 = v_CIN_2373_out0[15:15];
assign v__2505_out0 = v_CIN_2358_out0[0:0];
assign v__2520_out0 = v_CIN_2373_out0[0:0];
assign v__3054_out0 = v_CIN_2358_out0[9:9];
assign v__3069_out0 = v_CIN_2373_out0[9:9];
assign v__3088_out0 = v_CIN_2358_out0[2:2];
assign v__3103_out0 = v_CIN_2373_out0[2:2];
assign v__3142_out0 = v_CIN_2358_out0[7:7];
assign v__3157_out0 = v_CIN_2373_out0[7:7];
assign v__3826_out0 = v_CIN_2358_out0[1:1];
assign v__3841_out0 = v_CIN_2373_out0[1:1];
assign v__3864_out0 = v_CIN_2358_out0[10:10];
assign v__3879_out0 = v_CIN_2373_out0[10:10];
assign v__6803_out0 = v_CIN_2358_out0[11:11];
assign v__6818_out0 = v_CIN_2373_out0[11:11];
assign v__7647_out0 = v_CIN_2358_out0[12:12];
assign v__7662_out0 = v_CIN_2373_out0[12:12];
assign v__8702_out0 = v_CIN_2358_out0[13:13];
assign v__8717_out0 = v_CIN_2373_out0[13:13];
assign v__8772_out0 = v_CIN_2358_out0[14:14];
assign v__8787_out0 = v_CIN_2373_out0[14:14];
assign v__10722_out0 = v_CIN_2358_out0[5:5];
assign v__10737_out0 = v_CIN_2373_out0[5:5];
assign v__13451_out0 = v_CIN_2358_out0[4:4];
assign v__13466_out0 = v_CIN_2373_out0[4:4];
assign v_RM_3399_out0 = v__7647_out0;
assign v_RM_3400_out0 = v__8772_out0;
assign v_RM_3402_out0 = v__10722_out0;
assign v_RM_3403_out0 = v__13451_out0;
assign v_RM_3404_out0 = v__8702_out0;
assign v_RM_3405_out0 = v__3054_out0;
assign v_RM_3406_out0 = v__3864_out0;
assign v_RM_3407_out0 = v__3826_out0;
assign v_RM_3408_out0 = v__2158_out0;
assign v_RM_3409_out0 = v__1776_out0;
assign v_RM_3410_out0 = v__3142_out0;
assign v_RM_3411_out0 = v__6803_out0;
assign v_RM_3412_out0 = v__471_out0;
assign v_RM_3413_out0 = v__3088_out0;
assign v_RM_3623_out0 = v__7662_out0;
assign v_RM_3624_out0 = v__8787_out0;
assign v_RM_3626_out0 = v__10737_out0;
assign v_RM_3627_out0 = v__13466_out0;
assign v_RM_3628_out0 = v__8717_out0;
assign v_RM_3629_out0 = v__3069_out0;
assign v_RM_3630_out0 = v__3879_out0;
assign v_RM_3631_out0 = v__3841_out0;
assign v_RM_3632_out0 = v__2173_out0;
assign v_RM_3633_out0 = v__1791_out0;
assign v_RM_3634_out0 = v__3157_out0;
assign v_RM_3635_out0 = v__6818_out0;
assign v_RM_3636_out0 = v__486_out0;
assign v_RM_3637_out0 = v__3103_out0;
assign v_CIN_9854_out0 = v__2197_out0;
assign v_CIN_10078_out0 = v__2211_out0;
assign v_RM_11406_out0 = v__2505_out0;
assign v_RM_11870_out0 = v__2520_out0;
assign v_RD_5959_out0 = v_CIN_9854_out0;
assign v_RD_6423_out0 = v_CIN_10078_out0;
assign v_G1_7821_out0 = ((v_RD_5966_out0 && !v_RM_11406_out0) || (!v_RD_5966_out0) && v_RM_11406_out0);
assign v_G1_8285_out0 = ((v_RD_6430_out0 && !v_RM_11870_out0) || (!v_RD_6430_out0) && v_RM_11870_out0);
assign v_RM_11394_out0 = v_RM_3399_out0;
assign v_RM_11396_out0 = v_RM_3400_out0;
assign v_RM_11400_out0 = v_RM_3402_out0;
assign v_RM_11402_out0 = v_RM_3403_out0;
assign v_RM_11404_out0 = v_RM_3404_out0;
assign v_RM_11407_out0 = v_RM_3405_out0;
assign v_RM_11409_out0 = v_RM_3406_out0;
assign v_RM_11411_out0 = v_RM_3407_out0;
assign v_RM_11413_out0 = v_RM_3408_out0;
assign v_RM_11415_out0 = v_RM_3409_out0;
assign v_RM_11417_out0 = v_RM_3410_out0;
assign v_RM_11419_out0 = v_RM_3411_out0;
assign v_RM_11421_out0 = v_RM_3412_out0;
assign v_RM_11423_out0 = v_RM_3413_out0;
assign v_RM_11858_out0 = v_RM_3623_out0;
assign v_RM_11860_out0 = v_RM_3624_out0;
assign v_RM_11864_out0 = v_RM_3626_out0;
assign v_RM_11866_out0 = v_RM_3627_out0;
assign v_RM_11868_out0 = v_RM_3628_out0;
assign v_RM_11871_out0 = v_RM_3629_out0;
assign v_RM_11873_out0 = v_RM_3630_out0;
assign v_RM_11875_out0 = v_RM_3631_out0;
assign v_RM_11877_out0 = v_RM_3632_out0;
assign v_RM_11879_out0 = v_RM_3633_out0;
assign v_RM_11881_out0 = v_RM_3634_out0;
assign v_RM_11883_out0 = v_RM_3635_out0;
assign v_RM_11885_out0 = v_RM_3636_out0;
assign v_RM_11887_out0 = v_RM_3637_out0;
assign v_G2_12357_out0 = v_RD_5966_out0 && v_RM_11406_out0;
assign v_G2_12821_out0 = v_RD_6430_out0 && v_RM_11870_out0;
assign v_CARRY_4966_out0 = v_G2_12357_out0;
assign v_CARRY_5430_out0 = v_G2_12821_out0;
assign v_G1_7809_out0 = ((v_RD_5954_out0 && !v_RM_11394_out0) || (!v_RD_5954_out0) && v_RM_11394_out0);
assign v_G1_7811_out0 = ((v_RD_5956_out0 && !v_RM_11396_out0) || (!v_RD_5956_out0) && v_RM_11396_out0);
assign v_G1_7815_out0 = ((v_RD_5960_out0 && !v_RM_11400_out0) || (!v_RD_5960_out0) && v_RM_11400_out0);
assign v_G1_7817_out0 = ((v_RD_5962_out0 && !v_RM_11402_out0) || (!v_RD_5962_out0) && v_RM_11402_out0);
assign v_G1_7819_out0 = ((v_RD_5964_out0 && !v_RM_11404_out0) || (!v_RD_5964_out0) && v_RM_11404_out0);
assign v_G1_7822_out0 = ((v_RD_5967_out0 && !v_RM_11407_out0) || (!v_RD_5967_out0) && v_RM_11407_out0);
assign v_G1_7824_out0 = ((v_RD_5969_out0 && !v_RM_11409_out0) || (!v_RD_5969_out0) && v_RM_11409_out0);
assign v_G1_7826_out0 = ((v_RD_5971_out0 && !v_RM_11411_out0) || (!v_RD_5971_out0) && v_RM_11411_out0);
assign v_G1_7828_out0 = ((v_RD_5973_out0 && !v_RM_11413_out0) || (!v_RD_5973_out0) && v_RM_11413_out0);
assign v_G1_7830_out0 = ((v_RD_5975_out0 && !v_RM_11415_out0) || (!v_RD_5975_out0) && v_RM_11415_out0);
assign v_G1_7832_out0 = ((v_RD_5977_out0 && !v_RM_11417_out0) || (!v_RD_5977_out0) && v_RM_11417_out0);
assign v_G1_7834_out0 = ((v_RD_5979_out0 && !v_RM_11419_out0) || (!v_RD_5979_out0) && v_RM_11419_out0);
assign v_G1_7836_out0 = ((v_RD_5981_out0 && !v_RM_11421_out0) || (!v_RD_5981_out0) && v_RM_11421_out0);
assign v_G1_7838_out0 = ((v_RD_5983_out0 && !v_RM_11423_out0) || (!v_RD_5983_out0) && v_RM_11423_out0);
assign v_G1_8273_out0 = ((v_RD_6418_out0 && !v_RM_11858_out0) || (!v_RD_6418_out0) && v_RM_11858_out0);
assign v_G1_8275_out0 = ((v_RD_6420_out0 && !v_RM_11860_out0) || (!v_RD_6420_out0) && v_RM_11860_out0);
assign v_G1_8279_out0 = ((v_RD_6424_out0 && !v_RM_11864_out0) || (!v_RD_6424_out0) && v_RM_11864_out0);
assign v_G1_8281_out0 = ((v_RD_6426_out0 && !v_RM_11866_out0) || (!v_RD_6426_out0) && v_RM_11866_out0);
assign v_G1_8283_out0 = ((v_RD_6428_out0 && !v_RM_11868_out0) || (!v_RD_6428_out0) && v_RM_11868_out0);
assign v_G1_8286_out0 = ((v_RD_6431_out0 && !v_RM_11871_out0) || (!v_RD_6431_out0) && v_RM_11871_out0);
assign v_G1_8288_out0 = ((v_RD_6433_out0 && !v_RM_11873_out0) || (!v_RD_6433_out0) && v_RM_11873_out0);
assign v_G1_8290_out0 = ((v_RD_6435_out0 && !v_RM_11875_out0) || (!v_RD_6435_out0) && v_RM_11875_out0);
assign v_G1_8292_out0 = ((v_RD_6437_out0 && !v_RM_11877_out0) || (!v_RD_6437_out0) && v_RM_11877_out0);
assign v_G1_8294_out0 = ((v_RD_6439_out0 && !v_RM_11879_out0) || (!v_RD_6439_out0) && v_RM_11879_out0);
assign v_G1_8296_out0 = ((v_RD_6441_out0 && !v_RM_11881_out0) || (!v_RD_6441_out0) && v_RM_11881_out0);
assign v_G1_8298_out0 = ((v_RD_6443_out0 && !v_RM_11883_out0) || (!v_RD_6443_out0) && v_RM_11883_out0);
assign v_G1_8300_out0 = ((v_RD_6445_out0 && !v_RM_11885_out0) || (!v_RD_6445_out0) && v_RM_11885_out0);
assign v_G1_8302_out0 = ((v_RD_6447_out0 && !v_RM_11887_out0) || (!v_RD_6447_out0) && v_RM_11887_out0);
assign v_S_8967_out0 = v_G1_7821_out0;
assign v_S_9431_out0 = v_G1_8285_out0;
assign v_G2_12345_out0 = v_RD_5954_out0 && v_RM_11394_out0;
assign v_G2_12347_out0 = v_RD_5956_out0 && v_RM_11396_out0;
assign v_G2_12351_out0 = v_RD_5960_out0 && v_RM_11400_out0;
assign v_G2_12353_out0 = v_RD_5962_out0 && v_RM_11402_out0;
assign v_G2_12355_out0 = v_RD_5964_out0 && v_RM_11404_out0;
assign v_G2_12358_out0 = v_RD_5967_out0 && v_RM_11407_out0;
assign v_G2_12360_out0 = v_RD_5969_out0 && v_RM_11409_out0;
assign v_G2_12362_out0 = v_RD_5971_out0 && v_RM_11411_out0;
assign v_G2_12364_out0 = v_RD_5973_out0 && v_RM_11413_out0;
assign v_G2_12366_out0 = v_RD_5975_out0 && v_RM_11415_out0;
assign v_G2_12368_out0 = v_RD_5977_out0 && v_RM_11417_out0;
assign v_G2_12370_out0 = v_RD_5979_out0 && v_RM_11419_out0;
assign v_G2_12372_out0 = v_RD_5981_out0 && v_RM_11421_out0;
assign v_G2_12374_out0 = v_RD_5983_out0 && v_RM_11423_out0;
assign v_G2_12809_out0 = v_RD_6418_out0 && v_RM_11858_out0;
assign v_G2_12811_out0 = v_RD_6420_out0 && v_RM_11860_out0;
assign v_G2_12815_out0 = v_RD_6424_out0 && v_RM_11864_out0;
assign v_G2_12817_out0 = v_RD_6426_out0 && v_RM_11866_out0;
assign v_G2_12819_out0 = v_RD_6428_out0 && v_RM_11868_out0;
assign v_G2_12822_out0 = v_RD_6431_out0 && v_RM_11871_out0;
assign v_G2_12824_out0 = v_RD_6433_out0 && v_RM_11873_out0;
assign v_G2_12826_out0 = v_RD_6435_out0 && v_RM_11875_out0;
assign v_G2_12828_out0 = v_RD_6437_out0 && v_RM_11877_out0;
assign v_G2_12830_out0 = v_RD_6439_out0 && v_RM_11879_out0;
assign v_G2_12832_out0 = v_RD_6441_out0 && v_RM_11881_out0;
assign v_G2_12834_out0 = v_RD_6443_out0 && v_RM_11883_out0;
assign v_G2_12836_out0 = v_RD_6445_out0 && v_RM_11885_out0;
assign v_G2_12838_out0 = v_RD_6447_out0 && v_RM_11887_out0;
assign v_S_4668_out0 = v_S_8967_out0;
assign v_S_4683_out0 = v_S_9431_out0;
assign v_CARRY_4954_out0 = v_G2_12345_out0;
assign v_CARRY_4956_out0 = v_G2_12347_out0;
assign v_CARRY_4960_out0 = v_G2_12351_out0;
assign v_CARRY_4962_out0 = v_G2_12353_out0;
assign v_CARRY_4964_out0 = v_G2_12355_out0;
assign v_CARRY_4967_out0 = v_G2_12358_out0;
assign v_CARRY_4969_out0 = v_G2_12360_out0;
assign v_CARRY_4971_out0 = v_G2_12362_out0;
assign v_CARRY_4973_out0 = v_G2_12364_out0;
assign v_CARRY_4975_out0 = v_G2_12366_out0;
assign v_CARRY_4977_out0 = v_G2_12368_out0;
assign v_CARRY_4979_out0 = v_G2_12370_out0;
assign v_CARRY_4981_out0 = v_G2_12372_out0;
assign v_CARRY_4983_out0 = v_G2_12374_out0;
assign v_CARRY_5418_out0 = v_G2_12809_out0;
assign v_CARRY_5420_out0 = v_G2_12811_out0;
assign v_CARRY_5424_out0 = v_G2_12815_out0;
assign v_CARRY_5426_out0 = v_G2_12817_out0;
assign v_CARRY_5428_out0 = v_G2_12819_out0;
assign v_CARRY_5431_out0 = v_G2_12822_out0;
assign v_CARRY_5433_out0 = v_G2_12824_out0;
assign v_CARRY_5435_out0 = v_G2_12826_out0;
assign v_CARRY_5437_out0 = v_G2_12828_out0;
assign v_CARRY_5439_out0 = v_G2_12830_out0;
assign v_CARRY_5441_out0 = v_G2_12832_out0;
assign v_CARRY_5443_out0 = v_G2_12834_out0;
assign v_CARRY_5445_out0 = v_G2_12836_out0;
assign v_CARRY_5447_out0 = v_G2_12838_out0;
assign v_S_8955_out0 = v_G1_7809_out0;
assign v_S_8957_out0 = v_G1_7811_out0;
assign v_S_8961_out0 = v_G1_7815_out0;
assign v_S_8963_out0 = v_G1_7817_out0;
assign v_S_8965_out0 = v_G1_7819_out0;
assign v_S_8968_out0 = v_G1_7822_out0;
assign v_S_8970_out0 = v_G1_7824_out0;
assign v_S_8972_out0 = v_G1_7826_out0;
assign v_S_8974_out0 = v_G1_7828_out0;
assign v_S_8976_out0 = v_G1_7830_out0;
assign v_S_8978_out0 = v_G1_7832_out0;
assign v_S_8980_out0 = v_G1_7834_out0;
assign v_S_8982_out0 = v_G1_7836_out0;
assign v_S_8984_out0 = v_G1_7838_out0;
assign v_S_9419_out0 = v_G1_8273_out0;
assign v_S_9421_out0 = v_G1_8275_out0;
assign v_S_9425_out0 = v_G1_8279_out0;
assign v_S_9427_out0 = v_G1_8281_out0;
assign v_S_9429_out0 = v_G1_8283_out0;
assign v_S_9432_out0 = v_G1_8286_out0;
assign v_S_9434_out0 = v_G1_8288_out0;
assign v_S_9436_out0 = v_G1_8290_out0;
assign v_S_9438_out0 = v_G1_8292_out0;
assign v_S_9440_out0 = v_G1_8294_out0;
assign v_S_9442_out0 = v_G1_8296_out0;
assign v_S_9444_out0 = v_G1_8298_out0;
assign v_S_9446_out0 = v_G1_8300_out0;
assign v_S_9448_out0 = v_G1_8302_out0;
assign v_CIN_9860_out0 = v_CARRY_4966_out0;
assign v_CIN_10084_out0 = v_CARRY_5430_out0;
assign v__2439_out0 = { v__2191_out0,v_S_4668_out0 };
assign v__2440_out0 = { v__2192_out0,v_S_4683_out0 };
assign v_RD_5972_out0 = v_CIN_9860_out0;
assign v_RD_6436_out0 = v_CIN_10084_out0;
assign v_RM_11395_out0 = v_S_8955_out0;
assign v_RM_11397_out0 = v_S_8957_out0;
assign v_RM_11401_out0 = v_S_8961_out0;
assign v_RM_11403_out0 = v_S_8963_out0;
assign v_RM_11405_out0 = v_S_8965_out0;
assign v_RM_11408_out0 = v_S_8968_out0;
assign v_RM_11410_out0 = v_S_8970_out0;
assign v_RM_11412_out0 = v_S_8972_out0;
assign v_RM_11414_out0 = v_S_8974_out0;
assign v_RM_11416_out0 = v_S_8976_out0;
assign v_RM_11418_out0 = v_S_8978_out0;
assign v_RM_11420_out0 = v_S_8980_out0;
assign v_RM_11422_out0 = v_S_8982_out0;
assign v_RM_11424_out0 = v_S_8984_out0;
assign v_RM_11859_out0 = v_S_9419_out0;
assign v_RM_11861_out0 = v_S_9421_out0;
assign v_RM_11865_out0 = v_S_9425_out0;
assign v_RM_11867_out0 = v_S_9427_out0;
assign v_RM_11869_out0 = v_S_9429_out0;
assign v_RM_11872_out0 = v_S_9432_out0;
assign v_RM_11874_out0 = v_S_9434_out0;
assign v_RM_11876_out0 = v_S_9436_out0;
assign v_RM_11878_out0 = v_S_9438_out0;
assign v_RM_11880_out0 = v_S_9440_out0;
assign v_RM_11882_out0 = v_S_9442_out0;
assign v_RM_11884_out0 = v_S_9444_out0;
assign v_RM_11886_out0 = v_S_9446_out0;
assign v_RM_11888_out0 = v_S_9448_out0;
assign v_G1_7827_out0 = ((v_RD_5972_out0 && !v_RM_11412_out0) || (!v_RD_5972_out0) && v_RM_11412_out0);
assign v_G1_8291_out0 = ((v_RD_6436_out0 && !v_RM_11876_out0) || (!v_RD_6436_out0) && v_RM_11876_out0);
assign v_G2_12363_out0 = v_RD_5972_out0 && v_RM_11412_out0;
assign v_G2_12827_out0 = v_RD_6436_out0 && v_RM_11876_out0;
assign v_CARRY_4972_out0 = v_G2_12363_out0;
assign v_CARRY_5436_out0 = v_G2_12827_out0;
assign v_S_8973_out0 = v_G1_7827_out0;
assign v_S_9437_out0 = v_G1_8291_out0;
assign v_S_1271_out0 = v_S_8973_out0;
assign v_S_1495_out0 = v_S_9437_out0;
assign v_G1_4047_out0 = v_CARRY_4972_out0 || v_CARRY_4971_out0;
assign v_G1_4271_out0 = v_CARRY_5436_out0 || v_CARRY_5435_out0;
assign v_COUT_739_out0 = v_G1_4047_out0;
assign v_COUT_963_out0 = v_G1_4271_out0;
assign v_CIN_9866_out0 = v_COUT_739_out0;
assign v_CIN_10090_out0 = v_COUT_963_out0;
assign v_RD_5984_out0 = v_CIN_9866_out0;
assign v_RD_6448_out0 = v_CIN_10090_out0;
assign v_G1_7839_out0 = ((v_RD_5984_out0 && !v_RM_11424_out0) || (!v_RD_5984_out0) && v_RM_11424_out0);
assign v_G1_8303_out0 = ((v_RD_6448_out0 && !v_RM_11888_out0) || (!v_RD_6448_out0) && v_RM_11888_out0);
assign v_G2_12375_out0 = v_RD_5984_out0 && v_RM_11424_out0;
assign v_G2_12839_out0 = v_RD_6448_out0 && v_RM_11888_out0;
assign v_CARRY_4984_out0 = v_G2_12375_out0;
assign v_CARRY_5448_out0 = v_G2_12839_out0;
assign v_S_8985_out0 = v_G1_7839_out0;
assign v_S_9449_out0 = v_G1_8303_out0;
assign v_S_1277_out0 = v_S_8985_out0;
assign v_S_1501_out0 = v_S_9449_out0;
assign v_G1_4053_out0 = v_CARRY_4984_out0 || v_CARRY_4983_out0;
assign v_G1_4277_out0 = v_CARRY_5448_out0 || v_CARRY_5447_out0;
assign v_COUT_745_out0 = v_G1_4053_out0;
assign v_COUT_969_out0 = v_G1_4277_out0;
assign v__4785_out0 = { v_S_1271_out0,v_S_1277_out0 };
assign v__4800_out0 = { v_S_1495_out0,v_S_1501_out0 };
assign v_CIN_9861_out0 = v_COUT_745_out0;
assign v_CIN_10085_out0 = v_COUT_969_out0;
assign v_RD_5974_out0 = v_CIN_9861_out0;
assign v_RD_6438_out0 = v_CIN_10085_out0;
assign v_G1_7829_out0 = ((v_RD_5974_out0 && !v_RM_11414_out0) || (!v_RD_5974_out0) && v_RM_11414_out0);
assign v_G1_8293_out0 = ((v_RD_6438_out0 && !v_RM_11878_out0) || (!v_RD_6438_out0) && v_RM_11878_out0);
assign v_G2_12365_out0 = v_RD_5974_out0 && v_RM_11414_out0;
assign v_G2_12829_out0 = v_RD_6438_out0 && v_RM_11878_out0;
assign v_CARRY_4974_out0 = v_G2_12365_out0;
assign v_CARRY_5438_out0 = v_G2_12829_out0;
assign v_S_8975_out0 = v_G1_7829_out0;
assign v_S_9439_out0 = v_G1_8293_out0;
assign v_S_1272_out0 = v_S_8975_out0;
assign v_S_1496_out0 = v_S_9439_out0;
assign v_G1_4048_out0 = v_CARRY_4974_out0 || v_CARRY_4973_out0;
assign v_G1_4272_out0 = v_CARRY_5438_out0 || v_CARRY_5437_out0;
assign v_COUT_740_out0 = v_G1_4048_out0;
assign v_COUT_964_out0 = v_G1_4272_out0;
assign v__2555_out0 = { v__4785_out0,v_S_1272_out0 };
assign v__2570_out0 = { v__4800_out0,v_S_1496_out0 };
assign v_CIN_9856_out0 = v_COUT_740_out0;
assign v_CIN_10080_out0 = v_COUT_964_out0;
assign v_RD_5963_out0 = v_CIN_9856_out0;
assign v_RD_6427_out0 = v_CIN_10080_out0;
assign v_G1_7818_out0 = ((v_RD_5963_out0 && !v_RM_11403_out0) || (!v_RD_5963_out0) && v_RM_11403_out0);
assign v_G1_8282_out0 = ((v_RD_6427_out0 && !v_RM_11867_out0) || (!v_RD_6427_out0) && v_RM_11867_out0);
assign v_G2_12354_out0 = v_RD_5963_out0 && v_RM_11403_out0;
assign v_G2_12818_out0 = v_RD_6427_out0 && v_RM_11867_out0;
assign v_CARRY_4963_out0 = v_G2_12354_out0;
assign v_CARRY_5427_out0 = v_G2_12818_out0;
assign v_S_8964_out0 = v_G1_7818_out0;
assign v_S_9428_out0 = v_G1_8282_out0;
assign v_S_1267_out0 = v_S_8964_out0;
assign v_S_1491_out0 = v_S_9428_out0;
assign v_G1_4043_out0 = v_CARRY_4963_out0 || v_CARRY_4962_out0;
assign v_G1_4267_out0 = v_CARRY_5427_out0 || v_CARRY_5426_out0;
assign v_COUT_735_out0 = v_G1_4043_out0;
assign v_COUT_959_out0 = v_G1_4267_out0;
assign v__7035_out0 = { v__2555_out0,v_S_1267_out0 };
assign v__7050_out0 = { v__2570_out0,v_S_1491_out0 };
assign v_CIN_9855_out0 = v_COUT_735_out0;
assign v_CIN_10079_out0 = v_COUT_959_out0;
assign v_RD_5961_out0 = v_CIN_9855_out0;
assign v_RD_6425_out0 = v_CIN_10079_out0;
assign v_G1_7816_out0 = ((v_RD_5961_out0 && !v_RM_11401_out0) || (!v_RD_5961_out0) && v_RM_11401_out0);
assign v_G1_8280_out0 = ((v_RD_6425_out0 && !v_RM_11865_out0) || (!v_RD_6425_out0) && v_RM_11865_out0);
assign v_G2_12352_out0 = v_RD_5961_out0 && v_RM_11401_out0;
assign v_G2_12816_out0 = v_RD_6425_out0 && v_RM_11865_out0;
assign v_CARRY_4961_out0 = v_G2_12352_out0;
assign v_CARRY_5425_out0 = v_G2_12816_out0;
assign v_S_8962_out0 = v_G1_7816_out0;
assign v_S_9426_out0 = v_G1_8280_out0;
assign v_S_1266_out0 = v_S_8962_out0;
assign v_S_1490_out0 = v_S_9426_out0;
assign v_G1_4042_out0 = v_CARRY_4961_out0 || v_CARRY_4960_out0;
assign v_G1_4266_out0 = v_CARRY_5425_out0 || v_CARRY_5424_out0;
assign v_COUT_734_out0 = v_G1_4042_out0;
assign v_COUT_958_out0 = v_G1_4266_out0;
assign v__13521_out0 = { v__7035_out0,v_S_1266_out0 };
assign v__13536_out0 = { v__7050_out0,v_S_1490_out0 };
assign v_CIN_9862_out0 = v_COUT_734_out0;
assign v_CIN_10086_out0 = v_COUT_958_out0;
assign v_RD_5976_out0 = v_CIN_9862_out0;
assign v_RD_6440_out0 = v_CIN_10086_out0;
assign v_G1_7831_out0 = ((v_RD_5976_out0 && !v_RM_11416_out0) || (!v_RD_5976_out0) && v_RM_11416_out0);
assign v_G1_8295_out0 = ((v_RD_6440_out0 && !v_RM_11880_out0) || (!v_RD_6440_out0) && v_RM_11880_out0);
assign v_G2_12367_out0 = v_RD_5976_out0 && v_RM_11416_out0;
assign v_G2_12831_out0 = v_RD_6440_out0 && v_RM_11880_out0;
assign v_CARRY_4976_out0 = v_G2_12367_out0;
assign v_CARRY_5440_out0 = v_G2_12831_out0;
assign v_S_8977_out0 = v_G1_7831_out0;
assign v_S_9441_out0 = v_G1_8295_out0;
assign v_S_1273_out0 = v_S_8977_out0;
assign v_S_1497_out0 = v_S_9441_out0;
assign v_G1_4049_out0 = v_CARRY_4976_out0 || v_CARRY_4975_out0;
assign v_G1_4273_out0 = v_CARRY_5440_out0 || v_CARRY_5439_out0;
assign v_COUT_741_out0 = v_G1_4049_out0;
assign v_COUT_965_out0 = v_G1_4273_out0;
assign v__3314_out0 = { v__13521_out0,v_S_1273_out0 };
assign v__3329_out0 = { v__13536_out0,v_S_1497_out0 };
assign v_CIN_9863_out0 = v_COUT_741_out0;
assign v_CIN_10087_out0 = v_COUT_965_out0;
assign v_RD_5978_out0 = v_CIN_9863_out0;
assign v_RD_6442_out0 = v_CIN_10087_out0;
assign v_G1_7833_out0 = ((v_RD_5978_out0 && !v_RM_11418_out0) || (!v_RD_5978_out0) && v_RM_11418_out0);
assign v_G1_8297_out0 = ((v_RD_6442_out0 && !v_RM_11882_out0) || (!v_RD_6442_out0) && v_RM_11882_out0);
assign v_G2_12369_out0 = v_RD_5978_out0 && v_RM_11418_out0;
assign v_G2_12833_out0 = v_RD_6442_out0 && v_RM_11882_out0;
assign v_CARRY_4978_out0 = v_G2_12369_out0;
assign v_CARRY_5442_out0 = v_G2_12833_out0;
assign v_S_8979_out0 = v_G1_7833_out0;
assign v_S_9443_out0 = v_G1_8297_out0;
assign v_S_1274_out0 = v_S_8979_out0;
assign v_S_1498_out0 = v_S_9443_out0;
assign v_G1_4050_out0 = v_CARRY_4978_out0 || v_CARRY_4977_out0;
assign v_G1_4274_out0 = v_CARRY_5442_out0 || v_CARRY_5441_out0;
assign v_COUT_742_out0 = v_G1_4050_out0;
assign v_COUT_966_out0 = v_G1_4274_out0;
assign v__7150_out0 = { v__3314_out0,v_S_1274_out0 };
assign v__7165_out0 = { v__3329_out0,v_S_1498_out0 };
assign v_CIN_9865_out0 = v_COUT_742_out0;
assign v_CIN_10089_out0 = v_COUT_966_out0;
assign v_RD_5982_out0 = v_CIN_9865_out0;
assign v_RD_6446_out0 = v_CIN_10089_out0;
assign v_G1_7837_out0 = ((v_RD_5982_out0 && !v_RM_11422_out0) || (!v_RD_5982_out0) && v_RM_11422_out0);
assign v_G1_8301_out0 = ((v_RD_6446_out0 && !v_RM_11886_out0) || (!v_RD_6446_out0) && v_RM_11886_out0);
assign v_G2_12373_out0 = v_RD_5982_out0 && v_RM_11422_out0;
assign v_G2_12837_out0 = v_RD_6446_out0 && v_RM_11886_out0;
assign v_CARRY_4982_out0 = v_G2_12373_out0;
assign v_CARRY_5446_out0 = v_G2_12837_out0;
assign v_S_8983_out0 = v_G1_7837_out0;
assign v_S_9447_out0 = v_G1_8301_out0;
assign v_S_1276_out0 = v_S_8983_out0;
assign v_S_1500_out0 = v_S_9447_out0;
assign v_G1_4052_out0 = v_CARRY_4982_out0 || v_CARRY_4981_out0;
assign v_G1_4276_out0 = v_CARRY_5446_out0 || v_CARRY_5445_out0;
assign v_COUT_744_out0 = v_G1_4052_out0;
assign v_COUT_968_out0 = v_G1_4276_out0;
assign v__4752_out0 = { v__7150_out0,v_S_1276_out0 };
assign v__4767_out0 = { v__7165_out0,v_S_1500_out0 };
assign v_CIN_9858_out0 = v_COUT_744_out0;
assign v_CIN_10082_out0 = v_COUT_968_out0;
assign v_RD_5968_out0 = v_CIN_9858_out0;
assign v_RD_6432_out0 = v_CIN_10082_out0;
assign v_G1_7823_out0 = ((v_RD_5968_out0 && !v_RM_11408_out0) || (!v_RD_5968_out0) && v_RM_11408_out0);
assign v_G1_8287_out0 = ((v_RD_6432_out0 && !v_RM_11872_out0) || (!v_RD_6432_out0) && v_RM_11872_out0);
assign v_G2_12359_out0 = v_RD_5968_out0 && v_RM_11408_out0;
assign v_G2_12823_out0 = v_RD_6432_out0 && v_RM_11872_out0;
assign v_CARRY_4968_out0 = v_G2_12359_out0;
assign v_CARRY_5432_out0 = v_G2_12823_out0;
assign v_S_8969_out0 = v_G1_7823_out0;
assign v_S_9433_out0 = v_G1_8287_out0;
assign v_S_1269_out0 = v_S_8969_out0;
assign v_S_1493_out0 = v_S_9433_out0;
assign v_G1_4045_out0 = v_CARRY_4968_out0 || v_CARRY_4967_out0;
assign v_G1_4269_out0 = v_CARRY_5432_out0 || v_CARRY_5431_out0;
assign v_COUT_737_out0 = v_G1_4045_out0;
assign v_COUT_961_out0 = v_G1_4269_out0;
assign v__6929_out0 = { v__4752_out0,v_S_1269_out0 };
assign v__6944_out0 = { v__4767_out0,v_S_1493_out0 };
assign v_CIN_9859_out0 = v_COUT_737_out0;
assign v_CIN_10083_out0 = v_COUT_961_out0;
assign v_RD_5970_out0 = v_CIN_9859_out0;
assign v_RD_6434_out0 = v_CIN_10083_out0;
assign v_G1_7825_out0 = ((v_RD_5970_out0 && !v_RM_11410_out0) || (!v_RD_5970_out0) && v_RM_11410_out0);
assign v_G1_8289_out0 = ((v_RD_6434_out0 && !v_RM_11874_out0) || (!v_RD_6434_out0) && v_RM_11874_out0);
assign v_G2_12361_out0 = v_RD_5970_out0 && v_RM_11410_out0;
assign v_G2_12825_out0 = v_RD_6434_out0 && v_RM_11874_out0;
assign v_CARRY_4970_out0 = v_G2_12361_out0;
assign v_CARRY_5434_out0 = v_G2_12825_out0;
assign v_S_8971_out0 = v_G1_7825_out0;
assign v_S_9435_out0 = v_G1_8289_out0;
assign v_S_1270_out0 = v_S_8971_out0;
assign v_S_1494_out0 = v_S_9435_out0;
assign v_G1_4046_out0 = v_CARRY_4970_out0 || v_CARRY_4969_out0;
assign v_G1_4270_out0 = v_CARRY_5434_out0 || v_CARRY_5433_out0;
assign v_COUT_738_out0 = v_G1_4046_out0;
assign v_COUT_962_out0 = v_G1_4270_out0;
assign v__5805_out0 = { v__6929_out0,v_S_1270_out0 };
assign v__5820_out0 = { v__6944_out0,v_S_1494_out0 };
assign v_CIN_9864_out0 = v_COUT_738_out0;
assign v_CIN_10088_out0 = v_COUT_962_out0;
assign v_RD_5980_out0 = v_CIN_9864_out0;
assign v_RD_6444_out0 = v_CIN_10088_out0;
assign v_G1_7835_out0 = ((v_RD_5980_out0 && !v_RM_11420_out0) || (!v_RD_5980_out0) && v_RM_11420_out0);
assign v_G1_8299_out0 = ((v_RD_6444_out0 && !v_RM_11884_out0) || (!v_RD_6444_out0) && v_RM_11884_out0);
assign v_G2_12371_out0 = v_RD_5980_out0 && v_RM_11420_out0;
assign v_G2_12835_out0 = v_RD_6444_out0 && v_RM_11884_out0;
assign v_CARRY_4980_out0 = v_G2_12371_out0;
assign v_CARRY_5444_out0 = v_G2_12835_out0;
assign v_S_8981_out0 = v_G1_7835_out0;
assign v_S_9445_out0 = v_G1_8299_out0;
assign v_S_1275_out0 = v_S_8981_out0;
assign v_S_1499_out0 = v_S_9445_out0;
assign v_G1_4051_out0 = v_CARRY_4980_out0 || v_CARRY_4979_out0;
assign v_G1_4275_out0 = v_CARRY_5444_out0 || v_CARRY_5443_out0;
assign v_COUT_743_out0 = v_G1_4051_out0;
assign v_COUT_967_out0 = v_G1_4275_out0;
assign v__2029_out0 = { v__5805_out0,v_S_1275_out0 };
assign v__2044_out0 = { v__5820_out0,v_S_1499_out0 };
assign v_CIN_9852_out0 = v_COUT_743_out0;
assign v_CIN_10076_out0 = v_COUT_967_out0;
assign v_RD_5955_out0 = v_CIN_9852_out0;
assign v_RD_6419_out0 = v_CIN_10076_out0;
assign v_G1_7810_out0 = ((v_RD_5955_out0 && !v_RM_11395_out0) || (!v_RD_5955_out0) && v_RM_11395_out0);
assign v_G1_8274_out0 = ((v_RD_6419_out0 && !v_RM_11859_out0) || (!v_RD_6419_out0) && v_RM_11859_out0);
assign v_G2_12346_out0 = v_RD_5955_out0 && v_RM_11395_out0;
assign v_G2_12810_out0 = v_RD_6419_out0 && v_RM_11859_out0;
assign v_CARRY_4955_out0 = v_G2_12346_out0;
assign v_CARRY_5419_out0 = v_G2_12810_out0;
assign v_S_8956_out0 = v_G1_7810_out0;
assign v_S_9420_out0 = v_G1_8274_out0;
assign v_S_1263_out0 = v_S_8956_out0;
assign v_S_1487_out0 = v_S_9420_out0;
assign v_G1_4039_out0 = v_CARRY_4955_out0 || v_CARRY_4954_out0;
assign v_G1_4263_out0 = v_CARRY_5419_out0 || v_CARRY_5418_out0;
assign v_COUT_731_out0 = v_G1_4039_out0;
assign v_COUT_955_out0 = v_G1_4263_out0;
assign v__2796_out0 = { v__2029_out0,v_S_1263_out0 };
assign v__2811_out0 = { v__2044_out0,v_S_1487_out0 };
assign v_CIN_9857_out0 = v_COUT_731_out0;
assign v_CIN_10081_out0 = v_COUT_955_out0;
assign v_RD_5965_out0 = v_CIN_9857_out0;
assign v_RD_6429_out0 = v_CIN_10081_out0;
assign v_G1_7820_out0 = ((v_RD_5965_out0 && !v_RM_11405_out0) || (!v_RD_5965_out0) && v_RM_11405_out0);
assign v_G1_8284_out0 = ((v_RD_6429_out0 && !v_RM_11869_out0) || (!v_RD_6429_out0) && v_RM_11869_out0);
assign v_G2_12356_out0 = v_RD_5965_out0 && v_RM_11405_out0;
assign v_G2_12820_out0 = v_RD_6429_out0 && v_RM_11869_out0;
assign v_CARRY_4965_out0 = v_G2_12356_out0;
assign v_CARRY_5429_out0 = v_G2_12820_out0;
assign v_S_8966_out0 = v_G1_7820_out0;
assign v_S_9430_out0 = v_G1_8284_out0;
assign v_S_1268_out0 = v_S_8966_out0;
assign v_S_1492_out0 = v_S_9430_out0;
assign v_G1_4044_out0 = v_CARRY_4965_out0 || v_CARRY_4964_out0;
assign v_G1_4268_out0 = v_CARRY_5429_out0 || v_CARRY_5428_out0;
assign v_COUT_736_out0 = v_G1_4044_out0;
assign v_COUT_960_out0 = v_G1_4268_out0;
assign v__1828_out0 = { v__2796_out0,v_S_1268_out0 };
assign v__1843_out0 = { v__2811_out0,v_S_1492_out0 };
assign v_CIN_9853_out0 = v_COUT_736_out0;
assign v_CIN_10077_out0 = v_COUT_960_out0;
assign v_RD_5957_out0 = v_CIN_9853_out0;
assign v_RD_6421_out0 = v_CIN_10077_out0;
assign v_G1_7812_out0 = ((v_RD_5957_out0 && !v_RM_11397_out0) || (!v_RD_5957_out0) && v_RM_11397_out0);
assign v_G1_8276_out0 = ((v_RD_6421_out0 && !v_RM_11861_out0) || (!v_RD_6421_out0) && v_RM_11861_out0);
assign v_G2_12348_out0 = v_RD_5957_out0 && v_RM_11397_out0;
assign v_G2_12812_out0 = v_RD_6421_out0 && v_RM_11861_out0;
assign v_CARRY_4957_out0 = v_G2_12348_out0;
assign v_CARRY_5421_out0 = v_G2_12812_out0;
assign v_S_8958_out0 = v_G1_7812_out0;
assign v_S_9422_out0 = v_G1_8276_out0;
assign v_S_1264_out0 = v_S_8958_out0;
assign v_S_1488_out0 = v_S_9422_out0;
assign v_G1_4040_out0 = v_CARRY_4957_out0 || v_CARRY_4956_out0;
assign v_G1_4264_out0 = v_CARRY_5421_out0 || v_CARRY_5420_out0;
assign v_COUT_732_out0 = v_G1_4040_out0;
assign v_COUT_956_out0 = v_G1_4264_out0;
assign v__4552_out0 = { v__1828_out0,v_S_1264_out0 };
assign v__4567_out0 = { v__1843_out0,v_S_1488_out0 };
assign v_RM_3401_out0 = v_COUT_732_out0;
assign v_RM_3625_out0 = v_COUT_956_out0;
assign v_RM_11398_out0 = v_RM_3401_out0;
assign v_RM_11862_out0 = v_RM_3625_out0;
assign v_G1_7813_out0 = ((v_RD_5958_out0 && !v_RM_11398_out0) || (!v_RD_5958_out0) && v_RM_11398_out0);
assign v_G1_8277_out0 = ((v_RD_6422_out0 && !v_RM_11862_out0) || (!v_RD_6422_out0) && v_RM_11862_out0);
assign v_G2_12349_out0 = v_RD_5958_out0 && v_RM_11398_out0;
assign v_G2_12813_out0 = v_RD_6422_out0 && v_RM_11862_out0;
assign v_CARRY_4958_out0 = v_G2_12349_out0;
assign v_CARRY_5422_out0 = v_G2_12813_out0;
assign v_S_8959_out0 = v_G1_7813_out0;
assign v_S_9423_out0 = v_G1_8277_out0;
assign v_RM_11399_out0 = v_S_8959_out0;
assign v_RM_11863_out0 = v_S_9423_out0;
assign v_G1_7814_out0 = ((v_RD_5959_out0 && !v_RM_11399_out0) || (!v_RD_5959_out0) && v_RM_11399_out0);
assign v_G1_8278_out0 = ((v_RD_6423_out0 && !v_RM_11863_out0) || (!v_RD_6423_out0) && v_RM_11863_out0);
assign v_G2_12350_out0 = v_RD_5959_out0 && v_RM_11399_out0;
assign v_G2_12814_out0 = v_RD_6423_out0 && v_RM_11863_out0;
assign v_CARRY_4959_out0 = v_G2_12350_out0;
assign v_CARRY_5423_out0 = v_G2_12814_out0;
assign v_S_8960_out0 = v_G1_7814_out0;
assign v_S_9424_out0 = v_G1_8278_out0;
assign v_S_1265_out0 = v_S_8960_out0;
assign v_S_1489_out0 = v_S_9424_out0;
assign v_G1_4041_out0 = v_CARRY_4959_out0 || v_CARRY_4958_out0;
assign v_G1_4265_out0 = v_CARRY_5423_out0 || v_CARRY_5422_out0;
assign v_COUT_733_out0 = v_G1_4041_out0;
assign v_COUT_957_out0 = v_G1_4265_out0;
assign v__10654_out0 = { v__4552_out0,v_S_1265_out0 };
assign v__10669_out0 = { v__4567_out0,v_S_1489_out0 };
assign v__10949_out0 = { v__10654_out0,v_COUT_733_out0 };
assign v__10964_out0 = { v__10669_out0,v_COUT_957_out0 };
assign v_COUT_10919_out0 = v__10949_out0;
assign v_COUT_10934_out0 = v__10964_out0;
assign v_CIN_2363_out0 = v_COUT_10919_out0;
assign v_CIN_2378_out0 = v_COUT_10934_out0;
assign v__476_out0 = v_CIN_2363_out0[8:8];
assign v__491_out0 = v_CIN_2378_out0[8:8];
assign v__1781_out0 = v_CIN_2363_out0[6:6];
assign v__1796_out0 = v_CIN_2378_out0[6:6];
assign v__2163_out0 = v_CIN_2363_out0[3:3];
assign v__2178_out0 = v_CIN_2378_out0[3:3];
assign v__2202_out0 = v_CIN_2363_out0[15:15];
assign v__2216_out0 = v_CIN_2378_out0[15:15];
assign v__2510_out0 = v_CIN_2363_out0[0:0];
assign v__2525_out0 = v_CIN_2378_out0[0:0];
assign v__3059_out0 = v_CIN_2363_out0[9:9];
assign v__3074_out0 = v_CIN_2378_out0[9:9];
assign v__3093_out0 = v_CIN_2363_out0[2:2];
assign v__3108_out0 = v_CIN_2378_out0[2:2];
assign v__3147_out0 = v_CIN_2363_out0[7:7];
assign v__3162_out0 = v_CIN_2378_out0[7:7];
assign v__3831_out0 = v_CIN_2363_out0[1:1];
assign v__3846_out0 = v_CIN_2378_out0[1:1];
assign v__3869_out0 = v_CIN_2363_out0[10:10];
assign v__3884_out0 = v_CIN_2378_out0[10:10];
assign v__6808_out0 = v_CIN_2363_out0[11:11];
assign v__6823_out0 = v_CIN_2378_out0[11:11];
assign v__7652_out0 = v_CIN_2363_out0[12:12];
assign v__7667_out0 = v_CIN_2378_out0[12:12];
assign v__8707_out0 = v_CIN_2363_out0[13:13];
assign v__8722_out0 = v_CIN_2378_out0[13:13];
assign v__8777_out0 = v_CIN_2363_out0[14:14];
assign v__8792_out0 = v_CIN_2378_out0[14:14];
assign v__10727_out0 = v_CIN_2363_out0[5:5];
assign v__10742_out0 = v_CIN_2378_out0[5:5];
assign v__13456_out0 = v_CIN_2363_out0[4:4];
assign v__13471_out0 = v_CIN_2378_out0[4:4];
assign v_RM_3474_out0 = v__7652_out0;
assign v_RM_3475_out0 = v__8777_out0;
assign v_RM_3477_out0 = v__10727_out0;
assign v_RM_3478_out0 = v__13456_out0;
assign v_RM_3479_out0 = v__8707_out0;
assign v_RM_3480_out0 = v__3059_out0;
assign v_RM_3481_out0 = v__3869_out0;
assign v_RM_3482_out0 = v__3831_out0;
assign v_RM_3483_out0 = v__2163_out0;
assign v_RM_3484_out0 = v__1781_out0;
assign v_RM_3485_out0 = v__3147_out0;
assign v_RM_3486_out0 = v__6808_out0;
assign v_RM_3487_out0 = v__476_out0;
assign v_RM_3488_out0 = v__3093_out0;
assign v_RM_3698_out0 = v__7667_out0;
assign v_RM_3699_out0 = v__8792_out0;
assign v_RM_3701_out0 = v__10742_out0;
assign v_RM_3702_out0 = v__13471_out0;
assign v_RM_3703_out0 = v__8722_out0;
assign v_RM_3704_out0 = v__3074_out0;
assign v_RM_3705_out0 = v__3884_out0;
assign v_RM_3706_out0 = v__3846_out0;
assign v_RM_3707_out0 = v__2178_out0;
assign v_RM_3708_out0 = v__1796_out0;
assign v_RM_3709_out0 = v__3162_out0;
assign v_RM_3710_out0 = v__6823_out0;
assign v_RM_3711_out0 = v__491_out0;
assign v_RM_3712_out0 = v__3108_out0;
assign v_CIN_9929_out0 = v__2202_out0;
assign v_CIN_10153_out0 = v__2216_out0;
assign v_RM_11561_out0 = v__2510_out0;
assign v_RM_12025_out0 = v__2525_out0;
assign v_RD_6114_out0 = v_CIN_9929_out0;
assign v_RD_6578_out0 = v_CIN_10153_out0;
assign v_G1_7976_out0 = ((v_RD_6121_out0 && !v_RM_11561_out0) || (!v_RD_6121_out0) && v_RM_11561_out0);
assign v_G1_8440_out0 = ((v_RD_6585_out0 && !v_RM_12025_out0) || (!v_RD_6585_out0) && v_RM_12025_out0);
assign v_RM_11549_out0 = v_RM_3474_out0;
assign v_RM_11551_out0 = v_RM_3475_out0;
assign v_RM_11555_out0 = v_RM_3477_out0;
assign v_RM_11557_out0 = v_RM_3478_out0;
assign v_RM_11559_out0 = v_RM_3479_out0;
assign v_RM_11562_out0 = v_RM_3480_out0;
assign v_RM_11564_out0 = v_RM_3481_out0;
assign v_RM_11566_out0 = v_RM_3482_out0;
assign v_RM_11568_out0 = v_RM_3483_out0;
assign v_RM_11570_out0 = v_RM_3484_out0;
assign v_RM_11572_out0 = v_RM_3485_out0;
assign v_RM_11574_out0 = v_RM_3486_out0;
assign v_RM_11576_out0 = v_RM_3487_out0;
assign v_RM_11578_out0 = v_RM_3488_out0;
assign v_RM_12013_out0 = v_RM_3698_out0;
assign v_RM_12015_out0 = v_RM_3699_out0;
assign v_RM_12019_out0 = v_RM_3701_out0;
assign v_RM_12021_out0 = v_RM_3702_out0;
assign v_RM_12023_out0 = v_RM_3703_out0;
assign v_RM_12026_out0 = v_RM_3704_out0;
assign v_RM_12028_out0 = v_RM_3705_out0;
assign v_RM_12030_out0 = v_RM_3706_out0;
assign v_RM_12032_out0 = v_RM_3707_out0;
assign v_RM_12034_out0 = v_RM_3708_out0;
assign v_RM_12036_out0 = v_RM_3709_out0;
assign v_RM_12038_out0 = v_RM_3710_out0;
assign v_RM_12040_out0 = v_RM_3711_out0;
assign v_RM_12042_out0 = v_RM_3712_out0;
assign v_G2_12512_out0 = v_RD_6121_out0 && v_RM_11561_out0;
assign v_G2_12976_out0 = v_RD_6585_out0 && v_RM_12025_out0;
assign v_CARRY_5121_out0 = v_G2_12512_out0;
assign v_CARRY_5585_out0 = v_G2_12976_out0;
assign v_G1_7964_out0 = ((v_RD_6109_out0 && !v_RM_11549_out0) || (!v_RD_6109_out0) && v_RM_11549_out0);
assign v_G1_7966_out0 = ((v_RD_6111_out0 && !v_RM_11551_out0) || (!v_RD_6111_out0) && v_RM_11551_out0);
assign v_G1_7970_out0 = ((v_RD_6115_out0 && !v_RM_11555_out0) || (!v_RD_6115_out0) && v_RM_11555_out0);
assign v_G1_7972_out0 = ((v_RD_6117_out0 && !v_RM_11557_out0) || (!v_RD_6117_out0) && v_RM_11557_out0);
assign v_G1_7974_out0 = ((v_RD_6119_out0 && !v_RM_11559_out0) || (!v_RD_6119_out0) && v_RM_11559_out0);
assign v_G1_7977_out0 = ((v_RD_6122_out0 && !v_RM_11562_out0) || (!v_RD_6122_out0) && v_RM_11562_out0);
assign v_G1_7979_out0 = ((v_RD_6124_out0 && !v_RM_11564_out0) || (!v_RD_6124_out0) && v_RM_11564_out0);
assign v_G1_7981_out0 = ((v_RD_6126_out0 && !v_RM_11566_out0) || (!v_RD_6126_out0) && v_RM_11566_out0);
assign v_G1_7983_out0 = ((v_RD_6128_out0 && !v_RM_11568_out0) || (!v_RD_6128_out0) && v_RM_11568_out0);
assign v_G1_7985_out0 = ((v_RD_6130_out0 && !v_RM_11570_out0) || (!v_RD_6130_out0) && v_RM_11570_out0);
assign v_G1_7987_out0 = ((v_RD_6132_out0 && !v_RM_11572_out0) || (!v_RD_6132_out0) && v_RM_11572_out0);
assign v_G1_7989_out0 = ((v_RD_6134_out0 && !v_RM_11574_out0) || (!v_RD_6134_out0) && v_RM_11574_out0);
assign v_G1_7991_out0 = ((v_RD_6136_out0 && !v_RM_11576_out0) || (!v_RD_6136_out0) && v_RM_11576_out0);
assign v_G1_7993_out0 = ((v_RD_6138_out0 && !v_RM_11578_out0) || (!v_RD_6138_out0) && v_RM_11578_out0);
assign v_G1_8428_out0 = ((v_RD_6573_out0 && !v_RM_12013_out0) || (!v_RD_6573_out0) && v_RM_12013_out0);
assign v_G1_8430_out0 = ((v_RD_6575_out0 && !v_RM_12015_out0) || (!v_RD_6575_out0) && v_RM_12015_out0);
assign v_G1_8434_out0 = ((v_RD_6579_out0 && !v_RM_12019_out0) || (!v_RD_6579_out0) && v_RM_12019_out0);
assign v_G1_8436_out0 = ((v_RD_6581_out0 && !v_RM_12021_out0) || (!v_RD_6581_out0) && v_RM_12021_out0);
assign v_G1_8438_out0 = ((v_RD_6583_out0 && !v_RM_12023_out0) || (!v_RD_6583_out0) && v_RM_12023_out0);
assign v_G1_8441_out0 = ((v_RD_6586_out0 && !v_RM_12026_out0) || (!v_RD_6586_out0) && v_RM_12026_out0);
assign v_G1_8443_out0 = ((v_RD_6588_out0 && !v_RM_12028_out0) || (!v_RD_6588_out0) && v_RM_12028_out0);
assign v_G1_8445_out0 = ((v_RD_6590_out0 && !v_RM_12030_out0) || (!v_RD_6590_out0) && v_RM_12030_out0);
assign v_G1_8447_out0 = ((v_RD_6592_out0 && !v_RM_12032_out0) || (!v_RD_6592_out0) && v_RM_12032_out0);
assign v_G1_8449_out0 = ((v_RD_6594_out0 && !v_RM_12034_out0) || (!v_RD_6594_out0) && v_RM_12034_out0);
assign v_G1_8451_out0 = ((v_RD_6596_out0 && !v_RM_12036_out0) || (!v_RD_6596_out0) && v_RM_12036_out0);
assign v_G1_8453_out0 = ((v_RD_6598_out0 && !v_RM_12038_out0) || (!v_RD_6598_out0) && v_RM_12038_out0);
assign v_G1_8455_out0 = ((v_RD_6600_out0 && !v_RM_12040_out0) || (!v_RD_6600_out0) && v_RM_12040_out0);
assign v_G1_8457_out0 = ((v_RD_6602_out0 && !v_RM_12042_out0) || (!v_RD_6602_out0) && v_RM_12042_out0);
assign v_S_9122_out0 = v_G1_7976_out0;
assign v_S_9586_out0 = v_G1_8440_out0;
assign v_G2_12500_out0 = v_RD_6109_out0 && v_RM_11549_out0;
assign v_G2_12502_out0 = v_RD_6111_out0 && v_RM_11551_out0;
assign v_G2_12506_out0 = v_RD_6115_out0 && v_RM_11555_out0;
assign v_G2_12508_out0 = v_RD_6117_out0 && v_RM_11557_out0;
assign v_G2_12510_out0 = v_RD_6119_out0 && v_RM_11559_out0;
assign v_G2_12513_out0 = v_RD_6122_out0 && v_RM_11562_out0;
assign v_G2_12515_out0 = v_RD_6124_out0 && v_RM_11564_out0;
assign v_G2_12517_out0 = v_RD_6126_out0 && v_RM_11566_out0;
assign v_G2_12519_out0 = v_RD_6128_out0 && v_RM_11568_out0;
assign v_G2_12521_out0 = v_RD_6130_out0 && v_RM_11570_out0;
assign v_G2_12523_out0 = v_RD_6132_out0 && v_RM_11572_out0;
assign v_G2_12525_out0 = v_RD_6134_out0 && v_RM_11574_out0;
assign v_G2_12527_out0 = v_RD_6136_out0 && v_RM_11576_out0;
assign v_G2_12529_out0 = v_RD_6138_out0 && v_RM_11578_out0;
assign v_G2_12964_out0 = v_RD_6573_out0 && v_RM_12013_out0;
assign v_G2_12966_out0 = v_RD_6575_out0 && v_RM_12015_out0;
assign v_G2_12970_out0 = v_RD_6579_out0 && v_RM_12019_out0;
assign v_G2_12972_out0 = v_RD_6581_out0 && v_RM_12021_out0;
assign v_G2_12974_out0 = v_RD_6583_out0 && v_RM_12023_out0;
assign v_G2_12977_out0 = v_RD_6586_out0 && v_RM_12026_out0;
assign v_G2_12979_out0 = v_RD_6588_out0 && v_RM_12028_out0;
assign v_G2_12981_out0 = v_RD_6590_out0 && v_RM_12030_out0;
assign v_G2_12983_out0 = v_RD_6592_out0 && v_RM_12032_out0;
assign v_G2_12985_out0 = v_RD_6594_out0 && v_RM_12034_out0;
assign v_G2_12987_out0 = v_RD_6596_out0 && v_RM_12036_out0;
assign v_G2_12989_out0 = v_RD_6598_out0 && v_RM_12038_out0;
assign v_G2_12991_out0 = v_RD_6600_out0 && v_RM_12040_out0;
assign v_G2_12993_out0 = v_RD_6602_out0 && v_RM_12042_out0;
assign v_S_4673_out0 = v_S_9122_out0;
assign v_S_4688_out0 = v_S_9586_out0;
assign v_CARRY_5109_out0 = v_G2_12500_out0;
assign v_CARRY_5111_out0 = v_G2_12502_out0;
assign v_CARRY_5115_out0 = v_G2_12506_out0;
assign v_CARRY_5117_out0 = v_G2_12508_out0;
assign v_CARRY_5119_out0 = v_G2_12510_out0;
assign v_CARRY_5122_out0 = v_G2_12513_out0;
assign v_CARRY_5124_out0 = v_G2_12515_out0;
assign v_CARRY_5126_out0 = v_G2_12517_out0;
assign v_CARRY_5128_out0 = v_G2_12519_out0;
assign v_CARRY_5130_out0 = v_G2_12521_out0;
assign v_CARRY_5132_out0 = v_G2_12523_out0;
assign v_CARRY_5134_out0 = v_G2_12525_out0;
assign v_CARRY_5136_out0 = v_G2_12527_out0;
assign v_CARRY_5138_out0 = v_G2_12529_out0;
assign v_CARRY_5573_out0 = v_G2_12964_out0;
assign v_CARRY_5575_out0 = v_G2_12966_out0;
assign v_CARRY_5579_out0 = v_G2_12970_out0;
assign v_CARRY_5581_out0 = v_G2_12972_out0;
assign v_CARRY_5583_out0 = v_G2_12974_out0;
assign v_CARRY_5586_out0 = v_G2_12977_out0;
assign v_CARRY_5588_out0 = v_G2_12979_out0;
assign v_CARRY_5590_out0 = v_G2_12981_out0;
assign v_CARRY_5592_out0 = v_G2_12983_out0;
assign v_CARRY_5594_out0 = v_G2_12985_out0;
assign v_CARRY_5596_out0 = v_G2_12987_out0;
assign v_CARRY_5598_out0 = v_G2_12989_out0;
assign v_CARRY_5600_out0 = v_G2_12991_out0;
assign v_CARRY_5602_out0 = v_G2_12993_out0;
assign v_S_9110_out0 = v_G1_7964_out0;
assign v_S_9112_out0 = v_G1_7966_out0;
assign v_S_9116_out0 = v_G1_7970_out0;
assign v_S_9118_out0 = v_G1_7972_out0;
assign v_S_9120_out0 = v_G1_7974_out0;
assign v_S_9123_out0 = v_G1_7977_out0;
assign v_S_9125_out0 = v_G1_7979_out0;
assign v_S_9127_out0 = v_G1_7981_out0;
assign v_S_9129_out0 = v_G1_7983_out0;
assign v_S_9131_out0 = v_G1_7985_out0;
assign v_S_9133_out0 = v_G1_7987_out0;
assign v_S_9135_out0 = v_G1_7989_out0;
assign v_S_9137_out0 = v_G1_7991_out0;
assign v_S_9139_out0 = v_G1_7993_out0;
assign v_S_9574_out0 = v_G1_8428_out0;
assign v_S_9576_out0 = v_G1_8430_out0;
assign v_S_9580_out0 = v_G1_8434_out0;
assign v_S_9582_out0 = v_G1_8436_out0;
assign v_S_9584_out0 = v_G1_8438_out0;
assign v_S_9587_out0 = v_G1_8441_out0;
assign v_S_9589_out0 = v_G1_8443_out0;
assign v_S_9591_out0 = v_G1_8445_out0;
assign v_S_9593_out0 = v_G1_8447_out0;
assign v_S_9595_out0 = v_G1_8449_out0;
assign v_S_9597_out0 = v_G1_8451_out0;
assign v_S_9599_out0 = v_G1_8453_out0;
assign v_S_9601_out0 = v_G1_8455_out0;
assign v_S_9603_out0 = v_G1_8457_out0;
assign v_CIN_9935_out0 = v_CARRY_5121_out0;
assign v_CIN_10159_out0 = v_CARRY_5585_out0;
assign v_RD_6127_out0 = v_CIN_9935_out0;
assign v_RD_6591_out0 = v_CIN_10159_out0;
assign v__9802_out0 = { v__2439_out0,v_S_4673_out0 };
assign v__9803_out0 = { v__2440_out0,v_S_4688_out0 };
assign v_RM_11550_out0 = v_S_9110_out0;
assign v_RM_11552_out0 = v_S_9112_out0;
assign v_RM_11556_out0 = v_S_9116_out0;
assign v_RM_11558_out0 = v_S_9118_out0;
assign v_RM_11560_out0 = v_S_9120_out0;
assign v_RM_11563_out0 = v_S_9123_out0;
assign v_RM_11565_out0 = v_S_9125_out0;
assign v_RM_11567_out0 = v_S_9127_out0;
assign v_RM_11569_out0 = v_S_9129_out0;
assign v_RM_11571_out0 = v_S_9131_out0;
assign v_RM_11573_out0 = v_S_9133_out0;
assign v_RM_11575_out0 = v_S_9135_out0;
assign v_RM_11577_out0 = v_S_9137_out0;
assign v_RM_11579_out0 = v_S_9139_out0;
assign v_RM_12014_out0 = v_S_9574_out0;
assign v_RM_12016_out0 = v_S_9576_out0;
assign v_RM_12020_out0 = v_S_9580_out0;
assign v_RM_12022_out0 = v_S_9582_out0;
assign v_RM_12024_out0 = v_S_9584_out0;
assign v_RM_12027_out0 = v_S_9587_out0;
assign v_RM_12029_out0 = v_S_9589_out0;
assign v_RM_12031_out0 = v_S_9591_out0;
assign v_RM_12033_out0 = v_S_9593_out0;
assign v_RM_12035_out0 = v_S_9595_out0;
assign v_RM_12037_out0 = v_S_9597_out0;
assign v_RM_12039_out0 = v_S_9599_out0;
assign v_RM_12041_out0 = v_S_9601_out0;
assign v_RM_12043_out0 = v_S_9603_out0;
assign v_G1_7982_out0 = ((v_RD_6127_out0 && !v_RM_11567_out0) || (!v_RD_6127_out0) && v_RM_11567_out0);
assign v_G1_8446_out0 = ((v_RD_6591_out0 && !v_RM_12031_out0) || (!v_RD_6591_out0) && v_RM_12031_out0);
assign v_G2_12518_out0 = v_RD_6127_out0 && v_RM_11567_out0;
assign v_G2_12982_out0 = v_RD_6591_out0 && v_RM_12031_out0;
assign v_CARRY_5127_out0 = v_G2_12518_out0;
assign v_CARRY_5591_out0 = v_G2_12982_out0;
assign v_S_9128_out0 = v_G1_7982_out0;
assign v_S_9592_out0 = v_G1_8446_out0;
assign v_S_1346_out0 = v_S_9128_out0;
assign v_S_1570_out0 = v_S_9592_out0;
assign v_G1_4122_out0 = v_CARRY_5127_out0 || v_CARRY_5126_out0;
assign v_G1_4346_out0 = v_CARRY_5591_out0 || v_CARRY_5590_out0;
assign v_COUT_814_out0 = v_G1_4122_out0;
assign v_COUT_1038_out0 = v_G1_4346_out0;
assign v_CIN_9941_out0 = v_COUT_814_out0;
assign v_CIN_10165_out0 = v_COUT_1038_out0;
assign v_RD_6139_out0 = v_CIN_9941_out0;
assign v_RD_6603_out0 = v_CIN_10165_out0;
assign v_G1_7994_out0 = ((v_RD_6139_out0 && !v_RM_11579_out0) || (!v_RD_6139_out0) && v_RM_11579_out0);
assign v_G1_8458_out0 = ((v_RD_6603_out0 && !v_RM_12043_out0) || (!v_RD_6603_out0) && v_RM_12043_out0);
assign v_G2_12530_out0 = v_RD_6139_out0 && v_RM_11579_out0;
assign v_G2_12994_out0 = v_RD_6603_out0 && v_RM_12043_out0;
assign v_CARRY_5139_out0 = v_G2_12530_out0;
assign v_CARRY_5603_out0 = v_G2_12994_out0;
assign v_S_9140_out0 = v_G1_7994_out0;
assign v_S_9604_out0 = v_G1_8458_out0;
assign v_S_1352_out0 = v_S_9140_out0;
assign v_S_1576_out0 = v_S_9604_out0;
assign v_G1_4128_out0 = v_CARRY_5139_out0 || v_CARRY_5138_out0;
assign v_G1_4352_out0 = v_CARRY_5603_out0 || v_CARRY_5602_out0;
assign v_COUT_820_out0 = v_G1_4128_out0;
assign v_COUT_1044_out0 = v_G1_4352_out0;
assign v__4790_out0 = { v_S_1346_out0,v_S_1352_out0 };
assign v__4805_out0 = { v_S_1570_out0,v_S_1576_out0 };
assign v_CIN_9936_out0 = v_COUT_820_out0;
assign v_CIN_10160_out0 = v_COUT_1044_out0;
assign v_RD_6129_out0 = v_CIN_9936_out0;
assign v_RD_6593_out0 = v_CIN_10160_out0;
assign v_G1_7984_out0 = ((v_RD_6129_out0 && !v_RM_11569_out0) || (!v_RD_6129_out0) && v_RM_11569_out0);
assign v_G1_8448_out0 = ((v_RD_6593_out0 && !v_RM_12033_out0) || (!v_RD_6593_out0) && v_RM_12033_out0);
assign v_G2_12520_out0 = v_RD_6129_out0 && v_RM_11569_out0;
assign v_G2_12984_out0 = v_RD_6593_out0 && v_RM_12033_out0;
assign v_CARRY_5129_out0 = v_G2_12520_out0;
assign v_CARRY_5593_out0 = v_G2_12984_out0;
assign v_S_9130_out0 = v_G1_7984_out0;
assign v_S_9594_out0 = v_G1_8448_out0;
assign v_S_1347_out0 = v_S_9130_out0;
assign v_S_1571_out0 = v_S_9594_out0;
assign v_G1_4123_out0 = v_CARRY_5129_out0 || v_CARRY_5128_out0;
assign v_G1_4347_out0 = v_CARRY_5593_out0 || v_CARRY_5592_out0;
assign v_COUT_815_out0 = v_G1_4123_out0;
assign v_COUT_1039_out0 = v_G1_4347_out0;
assign v__2560_out0 = { v__4790_out0,v_S_1347_out0 };
assign v__2575_out0 = { v__4805_out0,v_S_1571_out0 };
assign v_CIN_9931_out0 = v_COUT_815_out0;
assign v_CIN_10155_out0 = v_COUT_1039_out0;
assign v_RD_6118_out0 = v_CIN_9931_out0;
assign v_RD_6582_out0 = v_CIN_10155_out0;
assign v_G1_7973_out0 = ((v_RD_6118_out0 && !v_RM_11558_out0) || (!v_RD_6118_out0) && v_RM_11558_out0);
assign v_G1_8437_out0 = ((v_RD_6582_out0 && !v_RM_12022_out0) || (!v_RD_6582_out0) && v_RM_12022_out0);
assign v_G2_12509_out0 = v_RD_6118_out0 && v_RM_11558_out0;
assign v_G2_12973_out0 = v_RD_6582_out0 && v_RM_12022_out0;
assign v_CARRY_5118_out0 = v_G2_12509_out0;
assign v_CARRY_5582_out0 = v_G2_12973_out0;
assign v_S_9119_out0 = v_G1_7973_out0;
assign v_S_9583_out0 = v_G1_8437_out0;
assign v_S_1342_out0 = v_S_9119_out0;
assign v_S_1566_out0 = v_S_9583_out0;
assign v_G1_4118_out0 = v_CARRY_5118_out0 || v_CARRY_5117_out0;
assign v_G1_4342_out0 = v_CARRY_5582_out0 || v_CARRY_5581_out0;
assign v_COUT_810_out0 = v_G1_4118_out0;
assign v_COUT_1034_out0 = v_G1_4342_out0;
assign v__7040_out0 = { v__2560_out0,v_S_1342_out0 };
assign v__7055_out0 = { v__2575_out0,v_S_1566_out0 };
assign v_CIN_9930_out0 = v_COUT_810_out0;
assign v_CIN_10154_out0 = v_COUT_1034_out0;
assign v_RD_6116_out0 = v_CIN_9930_out0;
assign v_RD_6580_out0 = v_CIN_10154_out0;
assign v_G1_7971_out0 = ((v_RD_6116_out0 && !v_RM_11556_out0) || (!v_RD_6116_out0) && v_RM_11556_out0);
assign v_G1_8435_out0 = ((v_RD_6580_out0 && !v_RM_12020_out0) || (!v_RD_6580_out0) && v_RM_12020_out0);
assign v_G2_12507_out0 = v_RD_6116_out0 && v_RM_11556_out0;
assign v_G2_12971_out0 = v_RD_6580_out0 && v_RM_12020_out0;
assign v_CARRY_5116_out0 = v_G2_12507_out0;
assign v_CARRY_5580_out0 = v_G2_12971_out0;
assign v_S_9117_out0 = v_G1_7971_out0;
assign v_S_9581_out0 = v_G1_8435_out0;
assign v_S_1341_out0 = v_S_9117_out0;
assign v_S_1565_out0 = v_S_9581_out0;
assign v_G1_4117_out0 = v_CARRY_5116_out0 || v_CARRY_5115_out0;
assign v_G1_4341_out0 = v_CARRY_5580_out0 || v_CARRY_5579_out0;
assign v_COUT_809_out0 = v_G1_4117_out0;
assign v_COUT_1033_out0 = v_G1_4341_out0;
assign v__13526_out0 = { v__7040_out0,v_S_1341_out0 };
assign v__13541_out0 = { v__7055_out0,v_S_1565_out0 };
assign v_CIN_9937_out0 = v_COUT_809_out0;
assign v_CIN_10161_out0 = v_COUT_1033_out0;
assign v_RD_6131_out0 = v_CIN_9937_out0;
assign v_RD_6595_out0 = v_CIN_10161_out0;
assign v_G1_7986_out0 = ((v_RD_6131_out0 && !v_RM_11571_out0) || (!v_RD_6131_out0) && v_RM_11571_out0);
assign v_G1_8450_out0 = ((v_RD_6595_out0 && !v_RM_12035_out0) || (!v_RD_6595_out0) && v_RM_12035_out0);
assign v_G2_12522_out0 = v_RD_6131_out0 && v_RM_11571_out0;
assign v_G2_12986_out0 = v_RD_6595_out0 && v_RM_12035_out0;
assign v_CARRY_5131_out0 = v_G2_12522_out0;
assign v_CARRY_5595_out0 = v_G2_12986_out0;
assign v_S_9132_out0 = v_G1_7986_out0;
assign v_S_9596_out0 = v_G1_8450_out0;
assign v_S_1348_out0 = v_S_9132_out0;
assign v_S_1572_out0 = v_S_9596_out0;
assign v_G1_4124_out0 = v_CARRY_5131_out0 || v_CARRY_5130_out0;
assign v_G1_4348_out0 = v_CARRY_5595_out0 || v_CARRY_5594_out0;
assign v_COUT_816_out0 = v_G1_4124_out0;
assign v_COUT_1040_out0 = v_G1_4348_out0;
assign v__3319_out0 = { v__13526_out0,v_S_1348_out0 };
assign v__3334_out0 = { v__13541_out0,v_S_1572_out0 };
assign v_CIN_9938_out0 = v_COUT_816_out0;
assign v_CIN_10162_out0 = v_COUT_1040_out0;
assign v_RD_6133_out0 = v_CIN_9938_out0;
assign v_RD_6597_out0 = v_CIN_10162_out0;
assign v_G1_7988_out0 = ((v_RD_6133_out0 && !v_RM_11573_out0) || (!v_RD_6133_out0) && v_RM_11573_out0);
assign v_G1_8452_out0 = ((v_RD_6597_out0 && !v_RM_12037_out0) || (!v_RD_6597_out0) && v_RM_12037_out0);
assign v_G2_12524_out0 = v_RD_6133_out0 && v_RM_11573_out0;
assign v_G2_12988_out0 = v_RD_6597_out0 && v_RM_12037_out0;
assign v_CARRY_5133_out0 = v_G2_12524_out0;
assign v_CARRY_5597_out0 = v_G2_12988_out0;
assign v_S_9134_out0 = v_G1_7988_out0;
assign v_S_9598_out0 = v_G1_8452_out0;
assign v_S_1349_out0 = v_S_9134_out0;
assign v_S_1573_out0 = v_S_9598_out0;
assign v_G1_4125_out0 = v_CARRY_5133_out0 || v_CARRY_5132_out0;
assign v_G1_4349_out0 = v_CARRY_5597_out0 || v_CARRY_5596_out0;
assign v_COUT_817_out0 = v_G1_4125_out0;
assign v_COUT_1041_out0 = v_G1_4349_out0;
assign v__7155_out0 = { v__3319_out0,v_S_1349_out0 };
assign v__7170_out0 = { v__3334_out0,v_S_1573_out0 };
assign v_CIN_9940_out0 = v_COUT_817_out0;
assign v_CIN_10164_out0 = v_COUT_1041_out0;
assign v_RD_6137_out0 = v_CIN_9940_out0;
assign v_RD_6601_out0 = v_CIN_10164_out0;
assign v_G1_7992_out0 = ((v_RD_6137_out0 && !v_RM_11577_out0) || (!v_RD_6137_out0) && v_RM_11577_out0);
assign v_G1_8456_out0 = ((v_RD_6601_out0 && !v_RM_12041_out0) || (!v_RD_6601_out0) && v_RM_12041_out0);
assign v_G2_12528_out0 = v_RD_6137_out0 && v_RM_11577_out0;
assign v_G2_12992_out0 = v_RD_6601_out0 && v_RM_12041_out0;
assign v_CARRY_5137_out0 = v_G2_12528_out0;
assign v_CARRY_5601_out0 = v_G2_12992_out0;
assign v_S_9138_out0 = v_G1_7992_out0;
assign v_S_9602_out0 = v_G1_8456_out0;
assign v_S_1351_out0 = v_S_9138_out0;
assign v_S_1575_out0 = v_S_9602_out0;
assign v_G1_4127_out0 = v_CARRY_5137_out0 || v_CARRY_5136_out0;
assign v_G1_4351_out0 = v_CARRY_5601_out0 || v_CARRY_5600_out0;
assign v_COUT_819_out0 = v_G1_4127_out0;
assign v_COUT_1043_out0 = v_G1_4351_out0;
assign v__4757_out0 = { v__7155_out0,v_S_1351_out0 };
assign v__4772_out0 = { v__7170_out0,v_S_1575_out0 };
assign v_CIN_9933_out0 = v_COUT_819_out0;
assign v_CIN_10157_out0 = v_COUT_1043_out0;
assign v_RD_6123_out0 = v_CIN_9933_out0;
assign v_RD_6587_out0 = v_CIN_10157_out0;
assign v_G1_7978_out0 = ((v_RD_6123_out0 && !v_RM_11563_out0) || (!v_RD_6123_out0) && v_RM_11563_out0);
assign v_G1_8442_out0 = ((v_RD_6587_out0 && !v_RM_12027_out0) || (!v_RD_6587_out0) && v_RM_12027_out0);
assign v_G2_12514_out0 = v_RD_6123_out0 && v_RM_11563_out0;
assign v_G2_12978_out0 = v_RD_6587_out0 && v_RM_12027_out0;
assign v_CARRY_5123_out0 = v_G2_12514_out0;
assign v_CARRY_5587_out0 = v_G2_12978_out0;
assign v_S_9124_out0 = v_G1_7978_out0;
assign v_S_9588_out0 = v_G1_8442_out0;
assign v_S_1344_out0 = v_S_9124_out0;
assign v_S_1568_out0 = v_S_9588_out0;
assign v_G1_4120_out0 = v_CARRY_5123_out0 || v_CARRY_5122_out0;
assign v_G1_4344_out0 = v_CARRY_5587_out0 || v_CARRY_5586_out0;
assign v_COUT_812_out0 = v_G1_4120_out0;
assign v_COUT_1036_out0 = v_G1_4344_out0;
assign v__6934_out0 = { v__4757_out0,v_S_1344_out0 };
assign v__6949_out0 = { v__4772_out0,v_S_1568_out0 };
assign v_CIN_9934_out0 = v_COUT_812_out0;
assign v_CIN_10158_out0 = v_COUT_1036_out0;
assign v_RD_6125_out0 = v_CIN_9934_out0;
assign v_RD_6589_out0 = v_CIN_10158_out0;
assign v_G1_7980_out0 = ((v_RD_6125_out0 && !v_RM_11565_out0) || (!v_RD_6125_out0) && v_RM_11565_out0);
assign v_G1_8444_out0 = ((v_RD_6589_out0 && !v_RM_12029_out0) || (!v_RD_6589_out0) && v_RM_12029_out0);
assign v_G2_12516_out0 = v_RD_6125_out0 && v_RM_11565_out0;
assign v_G2_12980_out0 = v_RD_6589_out0 && v_RM_12029_out0;
assign v_CARRY_5125_out0 = v_G2_12516_out0;
assign v_CARRY_5589_out0 = v_G2_12980_out0;
assign v_S_9126_out0 = v_G1_7980_out0;
assign v_S_9590_out0 = v_G1_8444_out0;
assign v_S_1345_out0 = v_S_9126_out0;
assign v_S_1569_out0 = v_S_9590_out0;
assign v_G1_4121_out0 = v_CARRY_5125_out0 || v_CARRY_5124_out0;
assign v_G1_4345_out0 = v_CARRY_5589_out0 || v_CARRY_5588_out0;
assign v_COUT_813_out0 = v_G1_4121_out0;
assign v_COUT_1037_out0 = v_G1_4345_out0;
assign v__5810_out0 = { v__6934_out0,v_S_1345_out0 };
assign v__5825_out0 = { v__6949_out0,v_S_1569_out0 };
assign v_CIN_9939_out0 = v_COUT_813_out0;
assign v_CIN_10163_out0 = v_COUT_1037_out0;
assign v_RD_6135_out0 = v_CIN_9939_out0;
assign v_RD_6599_out0 = v_CIN_10163_out0;
assign v_G1_7990_out0 = ((v_RD_6135_out0 && !v_RM_11575_out0) || (!v_RD_6135_out0) && v_RM_11575_out0);
assign v_G1_8454_out0 = ((v_RD_6599_out0 && !v_RM_12039_out0) || (!v_RD_6599_out0) && v_RM_12039_out0);
assign v_G2_12526_out0 = v_RD_6135_out0 && v_RM_11575_out0;
assign v_G2_12990_out0 = v_RD_6599_out0 && v_RM_12039_out0;
assign v_CARRY_5135_out0 = v_G2_12526_out0;
assign v_CARRY_5599_out0 = v_G2_12990_out0;
assign v_S_9136_out0 = v_G1_7990_out0;
assign v_S_9600_out0 = v_G1_8454_out0;
assign v_S_1350_out0 = v_S_9136_out0;
assign v_S_1574_out0 = v_S_9600_out0;
assign v_G1_4126_out0 = v_CARRY_5135_out0 || v_CARRY_5134_out0;
assign v_G1_4350_out0 = v_CARRY_5599_out0 || v_CARRY_5598_out0;
assign v_COUT_818_out0 = v_G1_4126_out0;
assign v_COUT_1042_out0 = v_G1_4350_out0;
assign v__2034_out0 = { v__5810_out0,v_S_1350_out0 };
assign v__2049_out0 = { v__5825_out0,v_S_1574_out0 };
assign v_CIN_9927_out0 = v_COUT_818_out0;
assign v_CIN_10151_out0 = v_COUT_1042_out0;
assign v_RD_6110_out0 = v_CIN_9927_out0;
assign v_RD_6574_out0 = v_CIN_10151_out0;
assign v_G1_7965_out0 = ((v_RD_6110_out0 && !v_RM_11550_out0) || (!v_RD_6110_out0) && v_RM_11550_out0);
assign v_G1_8429_out0 = ((v_RD_6574_out0 && !v_RM_12014_out0) || (!v_RD_6574_out0) && v_RM_12014_out0);
assign v_G2_12501_out0 = v_RD_6110_out0 && v_RM_11550_out0;
assign v_G2_12965_out0 = v_RD_6574_out0 && v_RM_12014_out0;
assign v_CARRY_5110_out0 = v_G2_12501_out0;
assign v_CARRY_5574_out0 = v_G2_12965_out0;
assign v_S_9111_out0 = v_G1_7965_out0;
assign v_S_9575_out0 = v_G1_8429_out0;
assign v_S_1338_out0 = v_S_9111_out0;
assign v_S_1562_out0 = v_S_9575_out0;
assign v_G1_4114_out0 = v_CARRY_5110_out0 || v_CARRY_5109_out0;
assign v_G1_4338_out0 = v_CARRY_5574_out0 || v_CARRY_5573_out0;
assign v_COUT_806_out0 = v_G1_4114_out0;
assign v_COUT_1030_out0 = v_G1_4338_out0;
assign v__2801_out0 = { v__2034_out0,v_S_1338_out0 };
assign v__2816_out0 = { v__2049_out0,v_S_1562_out0 };
assign v_CIN_9932_out0 = v_COUT_806_out0;
assign v_CIN_10156_out0 = v_COUT_1030_out0;
assign v_RD_6120_out0 = v_CIN_9932_out0;
assign v_RD_6584_out0 = v_CIN_10156_out0;
assign v_G1_7975_out0 = ((v_RD_6120_out0 && !v_RM_11560_out0) || (!v_RD_6120_out0) && v_RM_11560_out0);
assign v_G1_8439_out0 = ((v_RD_6584_out0 && !v_RM_12024_out0) || (!v_RD_6584_out0) && v_RM_12024_out0);
assign v_G2_12511_out0 = v_RD_6120_out0 && v_RM_11560_out0;
assign v_G2_12975_out0 = v_RD_6584_out0 && v_RM_12024_out0;
assign v_CARRY_5120_out0 = v_G2_12511_out0;
assign v_CARRY_5584_out0 = v_G2_12975_out0;
assign v_S_9121_out0 = v_G1_7975_out0;
assign v_S_9585_out0 = v_G1_8439_out0;
assign v_S_1343_out0 = v_S_9121_out0;
assign v_S_1567_out0 = v_S_9585_out0;
assign v_G1_4119_out0 = v_CARRY_5120_out0 || v_CARRY_5119_out0;
assign v_G1_4343_out0 = v_CARRY_5584_out0 || v_CARRY_5583_out0;
assign v_COUT_811_out0 = v_G1_4119_out0;
assign v_COUT_1035_out0 = v_G1_4343_out0;
assign v__1833_out0 = { v__2801_out0,v_S_1343_out0 };
assign v__1848_out0 = { v__2816_out0,v_S_1567_out0 };
assign v_CIN_9928_out0 = v_COUT_811_out0;
assign v_CIN_10152_out0 = v_COUT_1035_out0;
assign v_RD_6112_out0 = v_CIN_9928_out0;
assign v_RD_6576_out0 = v_CIN_10152_out0;
assign v_G1_7967_out0 = ((v_RD_6112_out0 && !v_RM_11552_out0) || (!v_RD_6112_out0) && v_RM_11552_out0);
assign v_G1_8431_out0 = ((v_RD_6576_out0 && !v_RM_12016_out0) || (!v_RD_6576_out0) && v_RM_12016_out0);
assign v_G2_12503_out0 = v_RD_6112_out0 && v_RM_11552_out0;
assign v_G2_12967_out0 = v_RD_6576_out0 && v_RM_12016_out0;
assign v_CARRY_5112_out0 = v_G2_12503_out0;
assign v_CARRY_5576_out0 = v_G2_12967_out0;
assign v_S_9113_out0 = v_G1_7967_out0;
assign v_S_9577_out0 = v_G1_8431_out0;
assign v_S_1339_out0 = v_S_9113_out0;
assign v_S_1563_out0 = v_S_9577_out0;
assign v_G1_4115_out0 = v_CARRY_5112_out0 || v_CARRY_5111_out0;
assign v_G1_4339_out0 = v_CARRY_5576_out0 || v_CARRY_5575_out0;
assign v_COUT_807_out0 = v_G1_4115_out0;
assign v_COUT_1031_out0 = v_G1_4339_out0;
assign v__4557_out0 = { v__1833_out0,v_S_1339_out0 };
assign v__4572_out0 = { v__1848_out0,v_S_1563_out0 };
assign v_RM_3476_out0 = v_COUT_807_out0;
assign v_RM_3700_out0 = v_COUT_1031_out0;
assign v_RM_11553_out0 = v_RM_3476_out0;
assign v_RM_12017_out0 = v_RM_3700_out0;
assign v_G1_7968_out0 = ((v_RD_6113_out0 && !v_RM_11553_out0) || (!v_RD_6113_out0) && v_RM_11553_out0);
assign v_G1_8432_out0 = ((v_RD_6577_out0 && !v_RM_12017_out0) || (!v_RD_6577_out0) && v_RM_12017_out0);
assign v_G2_12504_out0 = v_RD_6113_out0 && v_RM_11553_out0;
assign v_G2_12968_out0 = v_RD_6577_out0 && v_RM_12017_out0;
assign v_CARRY_5113_out0 = v_G2_12504_out0;
assign v_CARRY_5577_out0 = v_G2_12968_out0;
assign v_S_9114_out0 = v_G1_7968_out0;
assign v_S_9578_out0 = v_G1_8432_out0;
assign v_RM_11554_out0 = v_S_9114_out0;
assign v_RM_12018_out0 = v_S_9578_out0;
assign v_G1_7969_out0 = ((v_RD_6114_out0 && !v_RM_11554_out0) || (!v_RD_6114_out0) && v_RM_11554_out0);
assign v_G1_8433_out0 = ((v_RD_6578_out0 && !v_RM_12018_out0) || (!v_RD_6578_out0) && v_RM_12018_out0);
assign v_G2_12505_out0 = v_RD_6114_out0 && v_RM_11554_out0;
assign v_G2_12969_out0 = v_RD_6578_out0 && v_RM_12018_out0;
assign v_CARRY_5114_out0 = v_G2_12505_out0;
assign v_CARRY_5578_out0 = v_G2_12969_out0;
assign v_S_9115_out0 = v_G1_7969_out0;
assign v_S_9579_out0 = v_G1_8433_out0;
assign v_S_1340_out0 = v_S_9115_out0;
assign v_S_1564_out0 = v_S_9579_out0;
assign v_G1_4116_out0 = v_CARRY_5114_out0 || v_CARRY_5113_out0;
assign v_G1_4340_out0 = v_CARRY_5578_out0 || v_CARRY_5577_out0;
assign v_COUT_808_out0 = v_G1_4116_out0;
assign v_COUT_1032_out0 = v_G1_4340_out0;
assign v__10659_out0 = { v__4557_out0,v_S_1340_out0 };
assign v__10674_out0 = { v__4572_out0,v_S_1564_out0 };
assign v__10954_out0 = { v__10659_out0,v_COUT_808_out0 };
assign v__10969_out0 = { v__10674_out0,v_COUT_1032_out0 };
assign v_COUT_10924_out0 = v__10954_out0;
assign v_COUT_10939_out0 = v__10969_out0;
assign v_CIN_2367_out0 = v_COUT_10924_out0;
assign v_CIN_2382_out0 = v_COUT_10939_out0;
assign v__480_out0 = v_CIN_2367_out0[8:8];
assign v__495_out0 = v_CIN_2382_out0[8:8];
assign v__1785_out0 = v_CIN_2367_out0[6:6];
assign v__1800_out0 = v_CIN_2382_out0[6:6];
assign v__2167_out0 = v_CIN_2367_out0[3:3];
assign v__2182_out0 = v_CIN_2382_out0[3:3];
assign v__2206_out0 = v_CIN_2367_out0[15:15];
assign v__2220_out0 = v_CIN_2382_out0[15:15];
assign v__2514_out0 = v_CIN_2367_out0[0:0];
assign v__2529_out0 = v_CIN_2382_out0[0:0];
assign v__3063_out0 = v_CIN_2367_out0[9:9];
assign v__3078_out0 = v_CIN_2382_out0[9:9];
assign v__3097_out0 = v_CIN_2367_out0[2:2];
assign v__3112_out0 = v_CIN_2382_out0[2:2];
assign v__3151_out0 = v_CIN_2367_out0[7:7];
assign v__3166_out0 = v_CIN_2382_out0[7:7];
assign v__3835_out0 = v_CIN_2367_out0[1:1];
assign v__3850_out0 = v_CIN_2382_out0[1:1];
assign v__3873_out0 = v_CIN_2367_out0[10:10];
assign v__3888_out0 = v_CIN_2382_out0[10:10];
assign v__6812_out0 = v_CIN_2367_out0[11:11];
assign v__6827_out0 = v_CIN_2382_out0[11:11];
assign v__7656_out0 = v_CIN_2367_out0[12:12];
assign v__7671_out0 = v_CIN_2382_out0[12:12];
assign v__8711_out0 = v_CIN_2367_out0[13:13];
assign v__8726_out0 = v_CIN_2382_out0[13:13];
assign v__8781_out0 = v_CIN_2367_out0[14:14];
assign v__8796_out0 = v_CIN_2382_out0[14:14];
assign v__10731_out0 = v_CIN_2367_out0[5:5];
assign v__10746_out0 = v_CIN_2382_out0[5:5];
assign v__13460_out0 = v_CIN_2367_out0[4:4];
assign v__13475_out0 = v_CIN_2382_out0[4:4];
assign v_RM_3534_out0 = v__7656_out0;
assign v_RM_3535_out0 = v__8781_out0;
assign v_RM_3537_out0 = v__10731_out0;
assign v_RM_3538_out0 = v__13460_out0;
assign v_RM_3539_out0 = v__8711_out0;
assign v_RM_3540_out0 = v__3063_out0;
assign v_RM_3541_out0 = v__3873_out0;
assign v_RM_3542_out0 = v__3835_out0;
assign v_RM_3543_out0 = v__2167_out0;
assign v_RM_3544_out0 = v__1785_out0;
assign v_RM_3545_out0 = v__3151_out0;
assign v_RM_3546_out0 = v__6812_out0;
assign v_RM_3547_out0 = v__480_out0;
assign v_RM_3548_out0 = v__3097_out0;
assign v_RM_3758_out0 = v__7671_out0;
assign v_RM_3759_out0 = v__8796_out0;
assign v_RM_3761_out0 = v__10746_out0;
assign v_RM_3762_out0 = v__13475_out0;
assign v_RM_3763_out0 = v__8726_out0;
assign v_RM_3764_out0 = v__3078_out0;
assign v_RM_3765_out0 = v__3888_out0;
assign v_RM_3766_out0 = v__3850_out0;
assign v_RM_3767_out0 = v__2182_out0;
assign v_RM_3768_out0 = v__1800_out0;
assign v_RM_3769_out0 = v__3166_out0;
assign v_RM_3770_out0 = v__6827_out0;
assign v_RM_3771_out0 = v__495_out0;
assign v_RM_3772_out0 = v__3112_out0;
assign v_CIN_9989_out0 = v__2206_out0;
assign v_CIN_10213_out0 = v__2220_out0;
assign v_RM_11685_out0 = v__2514_out0;
assign v_RM_12149_out0 = v__2529_out0;
assign v_RD_6238_out0 = v_CIN_9989_out0;
assign v_RD_6702_out0 = v_CIN_10213_out0;
assign v_G1_8100_out0 = ((v_RD_6245_out0 && !v_RM_11685_out0) || (!v_RD_6245_out0) && v_RM_11685_out0);
assign v_G1_8564_out0 = ((v_RD_6709_out0 && !v_RM_12149_out0) || (!v_RD_6709_out0) && v_RM_12149_out0);
assign v_RM_11673_out0 = v_RM_3534_out0;
assign v_RM_11675_out0 = v_RM_3535_out0;
assign v_RM_11679_out0 = v_RM_3537_out0;
assign v_RM_11681_out0 = v_RM_3538_out0;
assign v_RM_11683_out0 = v_RM_3539_out0;
assign v_RM_11686_out0 = v_RM_3540_out0;
assign v_RM_11688_out0 = v_RM_3541_out0;
assign v_RM_11690_out0 = v_RM_3542_out0;
assign v_RM_11692_out0 = v_RM_3543_out0;
assign v_RM_11694_out0 = v_RM_3544_out0;
assign v_RM_11696_out0 = v_RM_3545_out0;
assign v_RM_11698_out0 = v_RM_3546_out0;
assign v_RM_11700_out0 = v_RM_3547_out0;
assign v_RM_11702_out0 = v_RM_3548_out0;
assign v_RM_12137_out0 = v_RM_3758_out0;
assign v_RM_12139_out0 = v_RM_3759_out0;
assign v_RM_12143_out0 = v_RM_3761_out0;
assign v_RM_12145_out0 = v_RM_3762_out0;
assign v_RM_12147_out0 = v_RM_3763_out0;
assign v_RM_12150_out0 = v_RM_3764_out0;
assign v_RM_12152_out0 = v_RM_3765_out0;
assign v_RM_12154_out0 = v_RM_3766_out0;
assign v_RM_12156_out0 = v_RM_3767_out0;
assign v_RM_12158_out0 = v_RM_3768_out0;
assign v_RM_12160_out0 = v_RM_3769_out0;
assign v_RM_12162_out0 = v_RM_3770_out0;
assign v_RM_12164_out0 = v_RM_3771_out0;
assign v_RM_12166_out0 = v_RM_3772_out0;
assign v_G2_12636_out0 = v_RD_6245_out0 && v_RM_11685_out0;
assign v_G2_13100_out0 = v_RD_6709_out0 && v_RM_12149_out0;
assign v_CARRY_5245_out0 = v_G2_12636_out0;
assign v_CARRY_5709_out0 = v_G2_13100_out0;
assign v_G1_8088_out0 = ((v_RD_6233_out0 && !v_RM_11673_out0) || (!v_RD_6233_out0) && v_RM_11673_out0);
assign v_G1_8090_out0 = ((v_RD_6235_out0 && !v_RM_11675_out0) || (!v_RD_6235_out0) && v_RM_11675_out0);
assign v_G1_8094_out0 = ((v_RD_6239_out0 && !v_RM_11679_out0) || (!v_RD_6239_out0) && v_RM_11679_out0);
assign v_G1_8096_out0 = ((v_RD_6241_out0 && !v_RM_11681_out0) || (!v_RD_6241_out0) && v_RM_11681_out0);
assign v_G1_8098_out0 = ((v_RD_6243_out0 && !v_RM_11683_out0) || (!v_RD_6243_out0) && v_RM_11683_out0);
assign v_G1_8101_out0 = ((v_RD_6246_out0 && !v_RM_11686_out0) || (!v_RD_6246_out0) && v_RM_11686_out0);
assign v_G1_8103_out0 = ((v_RD_6248_out0 && !v_RM_11688_out0) || (!v_RD_6248_out0) && v_RM_11688_out0);
assign v_G1_8105_out0 = ((v_RD_6250_out0 && !v_RM_11690_out0) || (!v_RD_6250_out0) && v_RM_11690_out0);
assign v_G1_8107_out0 = ((v_RD_6252_out0 && !v_RM_11692_out0) || (!v_RD_6252_out0) && v_RM_11692_out0);
assign v_G1_8109_out0 = ((v_RD_6254_out0 && !v_RM_11694_out0) || (!v_RD_6254_out0) && v_RM_11694_out0);
assign v_G1_8111_out0 = ((v_RD_6256_out0 && !v_RM_11696_out0) || (!v_RD_6256_out0) && v_RM_11696_out0);
assign v_G1_8113_out0 = ((v_RD_6258_out0 && !v_RM_11698_out0) || (!v_RD_6258_out0) && v_RM_11698_out0);
assign v_G1_8115_out0 = ((v_RD_6260_out0 && !v_RM_11700_out0) || (!v_RD_6260_out0) && v_RM_11700_out0);
assign v_G1_8117_out0 = ((v_RD_6262_out0 && !v_RM_11702_out0) || (!v_RD_6262_out0) && v_RM_11702_out0);
assign v_G1_8552_out0 = ((v_RD_6697_out0 && !v_RM_12137_out0) || (!v_RD_6697_out0) && v_RM_12137_out0);
assign v_G1_8554_out0 = ((v_RD_6699_out0 && !v_RM_12139_out0) || (!v_RD_6699_out0) && v_RM_12139_out0);
assign v_G1_8558_out0 = ((v_RD_6703_out0 && !v_RM_12143_out0) || (!v_RD_6703_out0) && v_RM_12143_out0);
assign v_G1_8560_out0 = ((v_RD_6705_out0 && !v_RM_12145_out0) || (!v_RD_6705_out0) && v_RM_12145_out0);
assign v_G1_8562_out0 = ((v_RD_6707_out0 && !v_RM_12147_out0) || (!v_RD_6707_out0) && v_RM_12147_out0);
assign v_G1_8565_out0 = ((v_RD_6710_out0 && !v_RM_12150_out0) || (!v_RD_6710_out0) && v_RM_12150_out0);
assign v_G1_8567_out0 = ((v_RD_6712_out0 && !v_RM_12152_out0) || (!v_RD_6712_out0) && v_RM_12152_out0);
assign v_G1_8569_out0 = ((v_RD_6714_out0 && !v_RM_12154_out0) || (!v_RD_6714_out0) && v_RM_12154_out0);
assign v_G1_8571_out0 = ((v_RD_6716_out0 && !v_RM_12156_out0) || (!v_RD_6716_out0) && v_RM_12156_out0);
assign v_G1_8573_out0 = ((v_RD_6718_out0 && !v_RM_12158_out0) || (!v_RD_6718_out0) && v_RM_12158_out0);
assign v_G1_8575_out0 = ((v_RD_6720_out0 && !v_RM_12160_out0) || (!v_RD_6720_out0) && v_RM_12160_out0);
assign v_G1_8577_out0 = ((v_RD_6722_out0 && !v_RM_12162_out0) || (!v_RD_6722_out0) && v_RM_12162_out0);
assign v_G1_8579_out0 = ((v_RD_6724_out0 && !v_RM_12164_out0) || (!v_RD_6724_out0) && v_RM_12164_out0);
assign v_G1_8581_out0 = ((v_RD_6726_out0 && !v_RM_12166_out0) || (!v_RD_6726_out0) && v_RM_12166_out0);
assign v_S_9246_out0 = v_G1_8100_out0;
assign v_S_9710_out0 = v_G1_8564_out0;
assign v_G2_12624_out0 = v_RD_6233_out0 && v_RM_11673_out0;
assign v_G2_12626_out0 = v_RD_6235_out0 && v_RM_11675_out0;
assign v_G2_12630_out0 = v_RD_6239_out0 && v_RM_11679_out0;
assign v_G2_12632_out0 = v_RD_6241_out0 && v_RM_11681_out0;
assign v_G2_12634_out0 = v_RD_6243_out0 && v_RM_11683_out0;
assign v_G2_12637_out0 = v_RD_6246_out0 && v_RM_11686_out0;
assign v_G2_12639_out0 = v_RD_6248_out0 && v_RM_11688_out0;
assign v_G2_12641_out0 = v_RD_6250_out0 && v_RM_11690_out0;
assign v_G2_12643_out0 = v_RD_6252_out0 && v_RM_11692_out0;
assign v_G2_12645_out0 = v_RD_6254_out0 && v_RM_11694_out0;
assign v_G2_12647_out0 = v_RD_6256_out0 && v_RM_11696_out0;
assign v_G2_12649_out0 = v_RD_6258_out0 && v_RM_11698_out0;
assign v_G2_12651_out0 = v_RD_6260_out0 && v_RM_11700_out0;
assign v_G2_12653_out0 = v_RD_6262_out0 && v_RM_11702_out0;
assign v_G2_13088_out0 = v_RD_6697_out0 && v_RM_12137_out0;
assign v_G2_13090_out0 = v_RD_6699_out0 && v_RM_12139_out0;
assign v_G2_13094_out0 = v_RD_6703_out0 && v_RM_12143_out0;
assign v_G2_13096_out0 = v_RD_6705_out0 && v_RM_12145_out0;
assign v_G2_13098_out0 = v_RD_6707_out0 && v_RM_12147_out0;
assign v_G2_13101_out0 = v_RD_6710_out0 && v_RM_12150_out0;
assign v_G2_13103_out0 = v_RD_6712_out0 && v_RM_12152_out0;
assign v_G2_13105_out0 = v_RD_6714_out0 && v_RM_12154_out0;
assign v_G2_13107_out0 = v_RD_6716_out0 && v_RM_12156_out0;
assign v_G2_13109_out0 = v_RD_6718_out0 && v_RM_12158_out0;
assign v_G2_13111_out0 = v_RD_6720_out0 && v_RM_12160_out0;
assign v_G2_13113_out0 = v_RD_6722_out0 && v_RM_12162_out0;
assign v_G2_13115_out0 = v_RD_6724_out0 && v_RM_12164_out0;
assign v_G2_13117_out0 = v_RD_6726_out0 && v_RM_12166_out0;
assign v_S_4677_out0 = v_S_9246_out0;
assign v_S_4692_out0 = v_S_9710_out0;
assign v_CARRY_5233_out0 = v_G2_12624_out0;
assign v_CARRY_5235_out0 = v_G2_12626_out0;
assign v_CARRY_5239_out0 = v_G2_12630_out0;
assign v_CARRY_5241_out0 = v_G2_12632_out0;
assign v_CARRY_5243_out0 = v_G2_12634_out0;
assign v_CARRY_5246_out0 = v_G2_12637_out0;
assign v_CARRY_5248_out0 = v_G2_12639_out0;
assign v_CARRY_5250_out0 = v_G2_12641_out0;
assign v_CARRY_5252_out0 = v_G2_12643_out0;
assign v_CARRY_5254_out0 = v_G2_12645_out0;
assign v_CARRY_5256_out0 = v_G2_12647_out0;
assign v_CARRY_5258_out0 = v_G2_12649_out0;
assign v_CARRY_5260_out0 = v_G2_12651_out0;
assign v_CARRY_5262_out0 = v_G2_12653_out0;
assign v_CARRY_5697_out0 = v_G2_13088_out0;
assign v_CARRY_5699_out0 = v_G2_13090_out0;
assign v_CARRY_5703_out0 = v_G2_13094_out0;
assign v_CARRY_5705_out0 = v_G2_13096_out0;
assign v_CARRY_5707_out0 = v_G2_13098_out0;
assign v_CARRY_5710_out0 = v_G2_13101_out0;
assign v_CARRY_5712_out0 = v_G2_13103_out0;
assign v_CARRY_5714_out0 = v_G2_13105_out0;
assign v_CARRY_5716_out0 = v_G2_13107_out0;
assign v_CARRY_5718_out0 = v_G2_13109_out0;
assign v_CARRY_5720_out0 = v_G2_13111_out0;
assign v_CARRY_5722_out0 = v_G2_13113_out0;
assign v_CARRY_5724_out0 = v_G2_13115_out0;
assign v_CARRY_5726_out0 = v_G2_13117_out0;
assign v_S_9234_out0 = v_G1_8088_out0;
assign v_S_9236_out0 = v_G1_8090_out0;
assign v_S_9240_out0 = v_G1_8094_out0;
assign v_S_9242_out0 = v_G1_8096_out0;
assign v_S_9244_out0 = v_G1_8098_out0;
assign v_S_9247_out0 = v_G1_8101_out0;
assign v_S_9249_out0 = v_G1_8103_out0;
assign v_S_9251_out0 = v_G1_8105_out0;
assign v_S_9253_out0 = v_G1_8107_out0;
assign v_S_9255_out0 = v_G1_8109_out0;
assign v_S_9257_out0 = v_G1_8111_out0;
assign v_S_9259_out0 = v_G1_8113_out0;
assign v_S_9261_out0 = v_G1_8115_out0;
assign v_S_9263_out0 = v_G1_8117_out0;
assign v_S_9698_out0 = v_G1_8552_out0;
assign v_S_9700_out0 = v_G1_8554_out0;
assign v_S_9704_out0 = v_G1_8558_out0;
assign v_S_9706_out0 = v_G1_8560_out0;
assign v_S_9708_out0 = v_G1_8562_out0;
assign v_S_9711_out0 = v_G1_8565_out0;
assign v_S_9713_out0 = v_G1_8567_out0;
assign v_S_9715_out0 = v_G1_8569_out0;
assign v_S_9717_out0 = v_G1_8571_out0;
assign v_S_9719_out0 = v_G1_8573_out0;
assign v_S_9721_out0 = v_G1_8575_out0;
assign v_S_9723_out0 = v_G1_8577_out0;
assign v_S_9725_out0 = v_G1_8579_out0;
assign v_S_9727_out0 = v_G1_8581_out0;
assign v_CIN_9995_out0 = v_CARRY_5245_out0;
assign v_CIN_10219_out0 = v_CARRY_5709_out0;
assign v_RD_6251_out0 = v_CIN_9995_out0;
assign v_RD_6715_out0 = v_CIN_10219_out0;
assign v__10767_out0 = { v__9802_out0,v_S_4677_out0 };
assign v__10768_out0 = { v__9803_out0,v_S_4692_out0 };
assign v_RM_11674_out0 = v_S_9234_out0;
assign v_RM_11676_out0 = v_S_9236_out0;
assign v_RM_11680_out0 = v_S_9240_out0;
assign v_RM_11682_out0 = v_S_9242_out0;
assign v_RM_11684_out0 = v_S_9244_out0;
assign v_RM_11687_out0 = v_S_9247_out0;
assign v_RM_11689_out0 = v_S_9249_out0;
assign v_RM_11691_out0 = v_S_9251_out0;
assign v_RM_11693_out0 = v_S_9253_out0;
assign v_RM_11695_out0 = v_S_9255_out0;
assign v_RM_11697_out0 = v_S_9257_out0;
assign v_RM_11699_out0 = v_S_9259_out0;
assign v_RM_11701_out0 = v_S_9261_out0;
assign v_RM_11703_out0 = v_S_9263_out0;
assign v_RM_12138_out0 = v_S_9698_out0;
assign v_RM_12140_out0 = v_S_9700_out0;
assign v_RM_12144_out0 = v_S_9704_out0;
assign v_RM_12146_out0 = v_S_9706_out0;
assign v_RM_12148_out0 = v_S_9708_out0;
assign v_RM_12151_out0 = v_S_9711_out0;
assign v_RM_12153_out0 = v_S_9713_out0;
assign v_RM_12155_out0 = v_S_9715_out0;
assign v_RM_12157_out0 = v_S_9717_out0;
assign v_RM_12159_out0 = v_S_9719_out0;
assign v_RM_12161_out0 = v_S_9721_out0;
assign v_RM_12163_out0 = v_S_9723_out0;
assign v_RM_12165_out0 = v_S_9725_out0;
assign v_RM_12167_out0 = v_S_9727_out0;
assign v_G1_8106_out0 = ((v_RD_6251_out0 && !v_RM_11691_out0) || (!v_RD_6251_out0) && v_RM_11691_out0);
assign v_G1_8570_out0 = ((v_RD_6715_out0 && !v_RM_12155_out0) || (!v_RD_6715_out0) && v_RM_12155_out0);
assign v_G2_12642_out0 = v_RD_6251_out0 && v_RM_11691_out0;
assign v_G2_13106_out0 = v_RD_6715_out0 && v_RM_12155_out0;
assign v_CARRY_5251_out0 = v_G2_12642_out0;
assign v_CARRY_5715_out0 = v_G2_13106_out0;
assign v_S_9252_out0 = v_G1_8106_out0;
assign v_S_9716_out0 = v_G1_8570_out0;
assign v_S_1406_out0 = v_S_9252_out0;
assign v_S_1630_out0 = v_S_9716_out0;
assign v_G1_4182_out0 = v_CARRY_5251_out0 || v_CARRY_5250_out0;
assign v_G1_4406_out0 = v_CARRY_5715_out0 || v_CARRY_5714_out0;
assign v_COUT_874_out0 = v_G1_4182_out0;
assign v_COUT_1098_out0 = v_G1_4406_out0;
assign v_CIN_10001_out0 = v_COUT_874_out0;
assign v_CIN_10225_out0 = v_COUT_1098_out0;
assign v_RD_6263_out0 = v_CIN_10001_out0;
assign v_RD_6727_out0 = v_CIN_10225_out0;
assign v_G1_8118_out0 = ((v_RD_6263_out0 && !v_RM_11703_out0) || (!v_RD_6263_out0) && v_RM_11703_out0);
assign v_G1_8582_out0 = ((v_RD_6727_out0 && !v_RM_12167_out0) || (!v_RD_6727_out0) && v_RM_12167_out0);
assign v_G2_12654_out0 = v_RD_6263_out0 && v_RM_11703_out0;
assign v_G2_13118_out0 = v_RD_6727_out0 && v_RM_12167_out0;
assign v_CARRY_5263_out0 = v_G2_12654_out0;
assign v_CARRY_5727_out0 = v_G2_13118_out0;
assign v_S_9264_out0 = v_G1_8118_out0;
assign v_S_9728_out0 = v_G1_8582_out0;
assign v_S_1412_out0 = v_S_9264_out0;
assign v_S_1636_out0 = v_S_9728_out0;
assign v_G1_4188_out0 = v_CARRY_5263_out0 || v_CARRY_5262_out0;
assign v_G1_4412_out0 = v_CARRY_5727_out0 || v_CARRY_5726_out0;
assign v_COUT_880_out0 = v_G1_4188_out0;
assign v_COUT_1104_out0 = v_G1_4412_out0;
assign v__4794_out0 = { v_S_1406_out0,v_S_1412_out0 };
assign v__4809_out0 = { v_S_1630_out0,v_S_1636_out0 };
assign v_CIN_9996_out0 = v_COUT_880_out0;
assign v_CIN_10220_out0 = v_COUT_1104_out0;
assign v_RD_6253_out0 = v_CIN_9996_out0;
assign v_RD_6717_out0 = v_CIN_10220_out0;
assign v_G1_8108_out0 = ((v_RD_6253_out0 && !v_RM_11693_out0) || (!v_RD_6253_out0) && v_RM_11693_out0);
assign v_G1_8572_out0 = ((v_RD_6717_out0 && !v_RM_12157_out0) || (!v_RD_6717_out0) && v_RM_12157_out0);
assign v_G2_12644_out0 = v_RD_6253_out0 && v_RM_11693_out0;
assign v_G2_13108_out0 = v_RD_6717_out0 && v_RM_12157_out0;
assign v_CARRY_5253_out0 = v_G2_12644_out0;
assign v_CARRY_5717_out0 = v_G2_13108_out0;
assign v_S_9254_out0 = v_G1_8108_out0;
assign v_S_9718_out0 = v_G1_8572_out0;
assign v_S_1407_out0 = v_S_9254_out0;
assign v_S_1631_out0 = v_S_9718_out0;
assign v_G1_4183_out0 = v_CARRY_5253_out0 || v_CARRY_5252_out0;
assign v_G1_4407_out0 = v_CARRY_5717_out0 || v_CARRY_5716_out0;
assign v_COUT_875_out0 = v_G1_4183_out0;
assign v_COUT_1099_out0 = v_G1_4407_out0;
assign v__2564_out0 = { v__4794_out0,v_S_1407_out0 };
assign v__2579_out0 = { v__4809_out0,v_S_1631_out0 };
assign v_CIN_9991_out0 = v_COUT_875_out0;
assign v_CIN_10215_out0 = v_COUT_1099_out0;
assign v_RD_6242_out0 = v_CIN_9991_out0;
assign v_RD_6706_out0 = v_CIN_10215_out0;
assign v_G1_8097_out0 = ((v_RD_6242_out0 && !v_RM_11682_out0) || (!v_RD_6242_out0) && v_RM_11682_out0);
assign v_G1_8561_out0 = ((v_RD_6706_out0 && !v_RM_12146_out0) || (!v_RD_6706_out0) && v_RM_12146_out0);
assign v_G2_12633_out0 = v_RD_6242_out0 && v_RM_11682_out0;
assign v_G2_13097_out0 = v_RD_6706_out0 && v_RM_12146_out0;
assign v_CARRY_5242_out0 = v_G2_12633_out0;
assign v_CARRY_5706_out0 = v_G2_13097_out0;
assign v_S_9243_out0 = v_G1_8097_out0;
assign v_S_9707_out0 = v_G1_8561_out0;
assign v_S_1402_out0 = v_S_9243_out0;
assign v_S_1626_out0 = v_S_9707_out0;
assign v_G1_4178_out0 = v_CARRY_5242_out0 || v_CARRY_5241_out0;
assign v_G1_4402_out0 = v_CARRY_5706_out0 || v_CARRY_5705_out0;
assign v_COUT_870_out0 = v_G1_4178_out0;
assign v_COUT_1094_out0 = v_G1_4402_out0;
assign v__7044_out0 = { v__2564_out0,v_S_1402_out0 };
assign v__7059_out0 = { v__2579_out0,v_S_1626_out0 };
assign v_CIN_9990_out0 = v_COUT_870_out0;
assign v_CIN_10214_out0 = v_COUT_1094_out0;
assign v_RD_6240_out0 = v_CIN_9990_out0;
assign v_RD_6704_out0 = v_CIN_10214_out0;
assign v_G1_8095_out0 = ((v_RD_6240_out0 && !v_RM_11680_out0) || (!v_RD_6240_out0) && v_RM_11680_out0);
assign v_G1_8559_out0 = ((v_RD_6704_out0 && !v_RM_12144_out0) || (!v_RD_6704_out0) && v_RM_12144_out0);
assign v_G2_12631_out0 = v_RD_6240_out0 && v_RM_11680_out0;
assign v_G2_13095_out0 = v_RD_6704_out0 && v_RM_12144_out0;
assign v_CARRY_5240_out0 = v_G2_12631_out0;
assign v_CARRY_5704_out0 = v_G2_13095_out0;
assign v_S_9241_out0 = v_G1_8095_out0;
assign v_S_9705_out0 = v_G1_8559_out0;
assign v_S_1401_out0 = v_S_9241_out0;
assign v_S_1625_out0 = v_S_9705_out0;
assign v_G1_4177_out0 = v_CARRY_5240_out0 || v_CARRY_5239_out0;
assign v_G1_4401_out0 = v_CARRY_5704_out0 || v_CARRY_5703_out0;
assign v_COUT_869_out0 = v_G1_4177_out0;
assign v_COUT_1093_out0 = v_G1_4401_out0;
assign v__13530_out0 = { v__7044_out0,v_S_1401_out0 };
assign v__13545_out0 = { v__7059_out0,v_S_1625_out0 };
assign v_CIN_9997_out0 = v_COUT_869_out0;
assign v_CIN_10221_out0 = v_COUT_1093_out0;
assign v_RD_6255_out0 = v_CIN_9997_out0;
assign v_RD_6719_out0 = v_CIN_10221_out0;
assign v_G1_8110_out0 = ((v_RD_6255_out0 && !v_RM_11695_out0) || (!v_RD_6255_out0) && v_RM_11695_out0);
assign v_G1_8574_out0 = ((v_RD_6719_out0 && !v_RM_12159_out0) || (!v_RD_6719_out0) && v_RM_12159_out0);
assign v_G2_12646_out0 = v_RD_6255_out0 && v_RM_11695_out0;
assign v_G2_13110_out0 = v_RD_6719_out0 && v_RM_12159_out0;
assign v_CARRY_5255_out0 = v_G2_12646_out0;
assign v_CARRY_5719_out0 = v_G2_13110_out0;
assign v_S_9256_out0 = v_G1_8110_out0;
assign v_S_9720_out0 = v_G1_8574_out0;
assign v_S_1408_out0 = v_S_9256_out0;
assign v_S_1632_out0 = v_S_9720_out0;
assign v_G1_4184_out0 = v_CARRY_5255_out0 || v_CARRY_5254_out0;
assign v_G1_4408_out0 = v_CARRY_5719_out0 || v_CARRY_5718_out0;
assign v_COUT_876_out0 = v_G1_4184_out0;
assign v_COUT_1100_out0 = v_G1_4408_out0;
assign v__3323_out0 = { v__13530_out0,v_S_1408_out0 };
assign v__3338_out0 = { v__13545_out0,v_S_1632_out0 };
assign v_CIN_9998_out0 = v_COUT_876_out0;
assign v_CIN_10222_out0 = v_COUT_1100_out0;
assign v_RD_6257_out0 = v_CIN_9998_out0;
assign v_RD_6721_out0 = v_CIN_10222_out0;
assign v_G1_8112_out0 = ((v_RD_6257_out0 && !v_RM_11697_out0) || (!v_RD_6257_out0) && v_RM_11697_out0);
assign v_G1_8576_out0 = ((v_RD_6721_out0 && !v_RM_12161_out0) || (!v_RD_6721_out0) && v_RM_12161_out0);
assign v_G2_12648_out0 = v_RD_6257_out0 && v_RM_11697_out0;
assign v_G2_13112_out0 = v_RD_6721_out0 && v_RM_12161_out0;
assign v_CARRY_5257_out0 = v_G2_12648_out0;
assign v_CARRY_5721_out0 = v_G2_13112_out0;
assign v_S_9258_out0 = v_G1_8112_out0;
assign v_S_9722_out0 = v_G1_8576_out0;
assign v_S_1409_out0 = v_S_9258_out0;
assign v_S_1633_out0 = v_S_9722_out0;
assign v_G1_4185_out0 = v_CARRY_5257_out0 || v_CARRY_5256_out0;
assign v_G1_4409_out0 = v_CARRY_5721_out0 || v_CARRY_5720_out0;
assign v_COUT_877_out0 = v_G1_4185_out0;
assign v_COUT_1101_out0 = v_G1_4409_out0;
assign v__7159_out0 = { v__3323_out0,v_S_1409_out0 };
assign v__7174_out0 = { v__3338_out0,v_S_1633_out0 };
assign v_CIN_10000_out0 = v_COUT_877_out0;
assign v_CIN_10224_out0 = v_COUT_1101_out0;
assign v_RD_6261_out0 = v_CIN_10000_out0;
assign v_RD_6725_out0 = v_CIN_10224_out0;
assign v_G1_8116_out0 = ((v_RD_6261_out0 && !v_RM_11701_out0) || (!v_RD_6261_out0) && v_RM_11701_out0);
assign v_G1_8580_out0 = ((v_RD_6725_out0 && !v_RM_12165_out0) || (!v_RD_6725_out0) && v_RM_12165_out0);
assign v_G2_12652_out0 = v_RD_6261_out0 && v_RM_11701_out0;
assign v_G2_13116_out0 = v_RD_6725_out0 && v_RM_12165_out0;
assign v_CARRY_5261_out0 = v_G2_12652_out0;
assign v_CARRY_5725_out0 = v_G2_13116_out0;
assign v_S_9262_out0 = v_G1_8116_out0;
assign v_S_9726_out0 = v_G1_8580_out0;
assign v_S_1411_out0 = v_S_9262_out0;
assign v_S_1635_out0 = v_S_9726_out0;
assign v_G1_4187_out0 = v_CARRY_5261_out0 || v_CARRY_5260_out0;
assign v_G1_4411_out0 = v_CARRY_5725_out0 || v_CARRY_5724_out0;
assign v_COUT_879_out0 = v_G1_4187_out0;
assign v_COUT_1103_out0 = v_G1_4411_out0;
assign v__4761_out0 = { v__7159_out0,v_S_1411_out0 };
assign v__4776_out0 = { v__7174_out0,v_S_1635_out0 };
assign v_CIN_9993_out0 = v_COUT_879_out0;
assign v_CIN_10217_out0 = v_COUT_1103_out0;
assign v_RD_6247_out0 = v_CIN_9993_out0;
assign v_RD_6711_out0 = v_CIN_10217_out0;
assign v_G1_8102_out0 = ((v_RD_6247_out0 && !v_RM_11687_out0) || (!v_RD_6247_out0) && v_RM_11687_out0);
assign v_G1_8566_out0 = ((v_RD_6711_out0 && !v_RM_12151_out0) || (!v_RD_6711_out0) && v_RM_12151_out0);
assign v_G2_12638_out0 = v_RD_6247_out0 && v_RM_11687_out0;
assign v_G2_13102_out0 = v_RD_6711_out0 && v_RM_12151_out0;
assign v_CARRY_5247_out0 = v_G2_12638_out0;
assign v_CARRY_5711_out0 = v_G2_13102_out0;
assign v_S_9248_out0 = v_G1_8102_out0;
assign v_S_9712_out0 = v_G1_8566_out0;
assign v_S_1404_out0 = v_S_9248_out0;
assign v_S_1628_out0 = v_S_9712_out0;
assign v_G1_4180_out0 = v_CARRY_5247_out0 || v_CARRY_5246_out0;
assign v_G1_4404_out0 = v_CARRY_5711_out0 || v_CARRY_5710_out0;
assign v_COUT_872_out0 = v_G1_4180_out0;
assign v_COUT_1096_out0 = v_G1_4404_out0;
assign v__6938_out0 = { v__4761_out0,v_S_1404_out0 };
assign v__6953_out0 = { v__4776_out0,v_S_1628_out0 };
assign v_CIN_9994_out0 = v_COUT_872_out0;
assign v_CIN_10218_out0 = v_COUT_1096_out0;
assign v_RD_6249_out0 = v_CIN_9994_out0;
assign v_RD_6713_out0 = v_CIN_10218_out0;
assign v_G1_8104_out0 = ((v_RD_6249_out0 && !v_RM_11689_out0) || (!v_RD_6249_out0) && v_RM_11689_out0);
assign v_G1_8568_out0 = ((v_RD_6713_out0 && !v_RM_12153_out0) || (!v_RD_6713_out0) && v_RM_12153_out0);
assign v_G2_12640_out0 = v_RD_6249_out0 && v_RM_11689_out0;
assign v_G2_13104_out0 = v_RD_6713_out0 && v_RM_12153_out0;
assign v_CARRY_5249_out0 = v_G2_12640_out0;
assign v_CARRY_5713_out0 = v_G2_13104_out0;
assign v_S_9250_out0 = v_G1_8104_out0;
assign v_S_9714_out0 = v_G1_8568_out0;
assign v_S_1405_out0 = v_S_9250_out0;
assign v_S_1629_out0 = v_S_9714_out0;
assign v_G1_4181_out0 = v_CARRY_5249_out0 || v_CARRY_5248_out0;
assign v_G1_4405_out0 = v_CARRY_5713_out0 || v_CARRY_5712_out0;
assign v_COUT_873_out0 = v_G1_4181_out0;
assign v_COUT_1097_out0 = v_G1_4405_out0;
assign v__5814_out0 = { v__6938_out0,v_S_1405_out0 };
assign v__5829_out0 = { v__6953_out0,v_S_1629_out0 };
assign v_CIN_9999_out0 = v_COUT_873_out0;
assign v_CIN_10223_out0 = v_COUT_1097_out0;
assign v_RD_6259_out0 = v_CIN_9999_out0;
assign v_RD_6723_out0 = v_CIN_10223_out0;
assign v_G1_8114_out0 = ((v_RD_6259_out0 && !v_RM_11699_out0) || (!v_RD_6259_out0) && v_RM_11699_out0);
assign v_G1_8578_out0 = ((v_RD_6723_out0 && !v_RM_12163_out0) || (!v_RD_6723_out0) && v_RM_12163_out0);
assign v_G2_12650_out0 = v_RD_6259_out0 && v_RM_11699_out0;
assign v_G2_13114_out0 = v_RD_6723_out0 && v_RM_12163_out0;
assign v_CARRY_5259_out0 = v_G2_12650_out0;
assign v_CARRY_5723_out0 = v_G2_13114_out0;
assign v_S_9260_out0 = v_G1_8114_out0;
assign v_S_9724_out0 = v_G1_8578_out0;
assign v_S_1410_out0 = v_S_9260_out0;
assign v_S_1634_out0 = v_S_9724_out0;
assign v_G1_4186_out0 = v_CARRY_5259_out0 || v_CARRY_5258_out0;
assign v_G1_4410_out0 = v_CARRY_5723_out0 || v_CARRY_5722_out0;
assign v_COUT_878_out0 = v_G1_4186_out0;
assign v_COUT_1102_out0 = v_G1_4410_out0;
assign v__2038_out0 = { v__5814_out0,v_S_1410_out0 };
assign v__2053_out0 = { v__5829_out0,v_S_1634_out0 };
assign v_CIN_9987_out0 = v_COUT_878_out0;
assign v_CIN_10211_out0 = v_COUT_1102_out0;
assign v_RD_6234_out0 = v_CIN_9987_out0;
assign v_RD_6698_out0 = v_CIN_10211_out0;
assign v_G1_8089_out0 = ((v_RD_6234_out0 && !v_RM_11674_out0) || (!v_RD_6234_out0) && v_RM_11674_out0);
assign v_G1_8553_out0 = ((v_RD_6698_out0 && !v_RM_12138_out0) || (!v_RD_6698_out0) && v_RM_12138_out0);
assign v_G2_12625_out0 = v_RD_6234_out0 && v_RM_11674_out0;
assign v_G2_13089_out0 = v_RD_6698_out0 && v_RM_12138_out0;
assign v_CARRY_5234_out0 = v_G2_12625_out0;
assign v_CARRY_5698_out0 = v_G2_13089_out0;
assign v_S_9235_out0 = v_G1_8089_out0;
assign v_S_9699_out0 = v_G1_8553_out0;
assign v_S_1398_out0 = v_S_9235_out0;
assign v_S_1622_out0 = v_S_9699_out0;
assign v_G1_4174_out0 = v_CARRY_5234_out0 || v_CARRY_5233_out0;
assign v_G1_4398_out0 = v_CARRY_5698_out0 || v_CARRY_5697_out0;
assign v_COUT_866_out0 = v_G1_4174_out0;
assign v_COUT_1090_out0 = v_G1_4398_out0;
assign v__2805_out0 = { v__2038_out0,v_S_1398_out0 };
assign v__2820_out0 = { v__2053_out0,v_S_1622_out0 };
assign v_CIN_9992_out0 = v_COUT_866_out0;
assign v_CIN_10216_out0 = v_COUT_1090_out0;
assign v_RD_6244_out0 = v_CIN_9992_out0;
assign v_RD_6708_out0 = v_CIN_10216_out0;
assign v_G1_8099_out0 = ((v_RD_6244_out0 && !v_RM_11684_out0) || (!v_RD_6244_out0) && v_RM_11684_out0);
assign v_G1_8563_out0 = ((v_RD_6708_out0 && !v_RM_12148_out0) || (!v_RD_6708_out0) && v_RM_12148_out0);
assign v_G2_12635_out0 = v_RD_6244_out0 && v_RM_11684_out0;
assign v_G2_13099_out0 = v_RD_6708_out0 && v_RM_12148_out0;
assign v_CARRY_5244_out0 = v_G2_12635_out0;
assign v_CARRY_5708_out0 = v_G2_13099_out0;
assign v_S_9245_out0 = v_G1_8099_out0;
assign v_S_9709_out0 = v_G1_8563_out0;
assign v_S_1403_out0 = v_S_9245_out0;
assign v_S_1627_out0 = v_S_9709_out0;
assign v_G1_4179_out0 = v_CARRY_5244_out0 || v_CARRY_5243_out0;
assign v_G1_4403_out0 = v_CARRY_5708_out0 || v_CARRY_5707_out0;
assign v_COUT_871_out0 = v_G1_4179_out0;
assign v_COUT_1095_out0 = v_G1_4403_out0;
assign v__1837_out0 = { v__2805_out0,v_S_1403_out0 };
assign v__1852_out0 = { v__2820_out0,v_S_1627_out0 };
assign v_CIN_9988_out0 = v_COUT_871_out0;
assign v_CIN_10212_out0 = v_COUT_1095_out0;
assign v_RD_6236_out0 = v_CIN_9988_out0;
assign v_RD_6700_out0 = v_CIN_10212_out0;
assign v_G1_8091_out0 = ((v_RD_6236_out0 && !v_RM_11676_out0) || (!v_RD_6236_out0) && v_RM_11676_out0);
assign v_G1_8555_out0 = ((v_RD_6700_out0 && !v_RM_12140_out0) || (!v_RD_6700_out0) && v_RM_12140_out0);
assign v_G2_12627_out0 = v_RD_6236_out0 && v_RM_11676_out0;
assign v_G2_13091_out0 = v_RD_6700_out0 && v_RM_12140_out0;
assign v_CARRY_5236_out0 = v_G2_12627_out0;
assign v_CARRY_5700_out0 = v_G2_13091_out0;
assign v_S_9237_out0 = v_G1_8091_out0;
assign v_S_9701_out0 = v_G1_8555_out0;
assign v_S_1399_out0 = v_S_9237_out0;
assign v_S_1623_out0 = v_S_9701_out0;
assign v_G1_4175_out0 = v_CARRY_5236_out0 || v_CARRY_5235_out0;
assign v_G1_4399_out0 = v_CARRY_5700_out0 || v_CARRY_5699_out0;
assign v_COUT_867_out0 = v_G1_4175_out0;
assign v_COUT_1091_out0 = v_G1_4399_out0;
assign v__4561_out0 = { v__1837_out0,v_S_1399_out0 };
assign v__4576_out0 = { v__1852_out0,v_S_1623_out0 };
assign v_RM_3536_out0 = v_COUT_867_out0;
assign v_RM_3760_out0 = v_COUT_1091_out0;
assign v_RM_11677_out0 = v_RM_3536_out0;
assign v_RM_12141_out0 = v_RM_3760_out0;
assign v_G1_8092_out0 = ((v_RD_6237_out0 && !v_RM_11677_out0) || (!v_RD_6237_out0) && v_RM_11677_out0);
assign v_G1_8556_out0 = ((v_RD_6701_out0 && !v_RM_12141_out0) || (!v_RD_6701_out0) && v_RM_12141_out0);
assign v_G2_12628_out0 = v_RD_6237_out0 && v_RM_11677_out0;
assign v_G2_13092_out0 = v_RD_6701_out0 && v_RM_12141_out0;
assign v_CARRY_5237_out0 = v_G2_12628_out0;
assign v_CARRY_5701_out0 = v_G2_13092_out0;
assign v_S_9238_out0 = v_G1_8092_out0;
assign v_S_9702_out0 = v_G1_8556_out0;
assign v_RM_11678_out0 = v_S_9238_out0;
assign v_RM_12142_out0 = v_S_9702_out0;
assign v_G1_8093_out0 = ((v_RD_6238_out0 && !v_RM_11678_out0) || (!v_RD_6238_out0) && v_RM_11678_out0);
assign v_G1_8557_out0 = ((v_RD_6702_out0 && !v_RM_12142_out0) || (!v_RD_6702_out0) && v_RM_12142_out0);
assign v_G2_12629_out0 = v_RD_6238_out0 && v_RM_11678_out0;
assign v_G2_13093_out0 = v_RD_6702_out0 && v_RM_12142_out0;
assign v_CARRY_5238_out0 = v_G2_12629_out0;
assign v_CARRY_5702_out0 = v_G2_13093_out0;
assign v_S_9239_out0 = v_G1_8093_out0;
assign v_S_9703_out0 = v_G1_8557_out0;
assign v_S_1400_out0 = v_S_9239_out0;
assign v_S_1624_out0 = v_S_9703_out0;
assign v_G1_4176_out0 = v_CARRY_5238_out0 || v_CARRY_5237_out0;
assign v_G1_4400_out0 = v_CARRY_5702_out0 || v_CARRY_5701_out0;
assign v_COUT_868_out0 = v_G1_4176_out0;
assign v_COUT_1092_out0 = v_G1_4400_out0;
assign v__10663_out0 = { v__4561_out0,v_S_1400_out0 };
assign v__10678_out0 = { v__4576_out0,v_S_1624_out0 };
assign v__10958_out0 = { v__10663_out0,v_COUT_868_out0 };
assign v__10973_out0 = { v__10678_out0,v_COUT_1092_out0 };
assign v_COUT_10928_out0 = v__10958_out0;
assign v_COUT_10943_out0 = v__10973_out0;
assign v_CIN_2362_out0 = v_COUT_10928_out0;
assign v_CIN_2377_out0 = v_COUT_10943_out0;
assign v__475_out0 = v_CIN_2362_out0[8:8];
assign v__490_out0 = v_CIN_2377_out0[8:8];
assign v__1780_out0 = v_CIN_2362_out0[6:6];
assign v__1795_out0 = v_CIN_2377_out0[6:6];
assign v__2162_out0 = v_CIN_2362_out0[3:3];
assign v__2177_out0 = v_CIN_2377_out0[3:3];
assign v__2201_out0 = v_CIN_2362_out0[15:15];
assign v__2215_out0 = v_CIN_2377_out0[15:15];
assign v__2509_out0 = v_CIN_2362_out0[0:0];
assign v__2524_out0 = v_CIN_2377_out0[0:0];
assign v__3058_out0 = v_CIN_2362_out0[9:9];
assign v__3073_out0 = v_CIN_2377_out0[9:9];
assign v__3092_out0 = v_CIN_2362_out0[2:2];
assign v__3107_out0 = v_CIN_2377_out0[2:2];
assign v__3146_out0 = v_CIN_2362_out0[7:7];
assign v__3161_out0 = v_CIN_2377_out0[7:7];
assign v__3830_out0 = v_CIN_2362_out0[1:1];
assign v__3845_out0 = v_CIN_2377_out0[1:1];
assign v__3868_out0 = v_CIN_2362_out0[10:10];
assign v__3883_out0 = v_CIN_2377_out0[10:10];
assign v__6807_out0 = v_CIN_2362_out0[11:11];
assign v__6822_out0 = v_CIN_2377_out0[11:11];
assign v__7651_out0 = v_CIN_2362_out0[12:12];
assign v__7666_out0 = v_CIN_2377_out0[12:12];
assign v__8706_out0 = v_CIN_2362_out0[13:13];
assign v__8721_out0 = v_CIN_2377_out0[13:13];
assign v__8776_out0 = v_CIN_2362_out0[14:14];
assign v__8791_out0 = v_CIN_2377_out0[14:14];
assign v__10726_out0 = v_CIN_2362_out0[5:5];
assign v__10741_out0 = v_CIN_2377_out0[5:5];
assign v__13455_out0 = v_CIN_2362_out0[4:4];
assign v__13470_out0 = v_CIN_2377_out0[4:4];
assign v_RM_3459_out0 = v__7651_out0;
assign v_RM_3460_out0 = v__8776_out0;
assign v_RM_3462_out0 = v__10726_out0;
assign v_RM_3463_out0 = v__13455_out0;
assign v_RM_3464_out0 = v__8706_out0;
assign v_RM_3465_out0 = v__3058_out0;
assign v_RM_3466_out0 = v__3868_out0;
assign v_RM_3467_out0 = v__3830_out0;
assign v_RM_3468_out0 = v__2162_out0;
assign v_RM_3469_out0 = v__1780_out0;
assign v_RM_3470_out0 = v__3146_out0;
assign v_RM_3471_out0 = v__6807_out0;
assign v_RM_3472_out0 = v__475_out0;
assign v_RM_3473_out0 = v__3092_out0;
assign v_RM_3683_out0 = v__7666_out0;
assign v_RM_3684_out0 = v__8791_out0;
assign v_RM_3686_out0 = v__10741_out0;
assign v_RM_3687_out0 = v__13470_out0;
assign v_RM_3688_out0 = v__8721_out0;
assign v_RM_3689_out0 = v__3073_out0;
assign v_RM_3690_out0 = v__3883_out0;
assign v_RM_3691_out0 = v__3845_out0;
assign v_RM_3692_out0 = v__2177_out0;
assign v_RM_3693_out0 = v__1795_out0;
assign v_RM_3694_out0 = v__3161_out0;
assign v_RM_3695_out0 = v__6822_out0;
assign v_RM_3696_out0 = v__490_out0;
assign v_RM_3697_out0 = v__3107_out0;
assign v_CIN_9914_out0 = v__2201_out0;
assign v_CIN_10138_out0 = v__2215_out0;
assign v_RM_11530_out0 = v__2509_out0;
assign v_RM_11994_out0 = v__2524_out0;
assign v_RD_6083_out0 = v_CIN_9914_out0;
assign v_RD_6547_out0 = v_CIN_10138_out0;
assign v_G1_7945_out0 = ((v_RD_6090_out0 && !v_RM_11530_out0) || (!v_RD_6090_out0) && v_RM_11530_out0);
assign v_G1_8409_out0 = ((v_RD_6554_out0 && !v_RM_11994_out0) || (!v_RD_6554_out0) && v_RM_11994_out0);
assign v_RM_11518_out0 = v_RM_3459_out0;
assign v_RM_11520_out0 = v_RM_3460_out0;
assign v_RM_11524_out0 = v_RM_3462_out0;
assign v_RM_11526_out0 = v_RM_3463_out0;
assign v_RM_11528_out0 = v_RM_3464_out0;
assign v_RM_11531_out0 = v_RM_3465_out0;
assign v_RM_11533_out0 = v_RM_3466_out0;
assign v_RM_11535_out0 = v_RM_3467_out0;
assign v_RM_11537_out0 = v_RM_3468_out0;
assign v_RM_11539_out0 = v_RM_3469_out0;
assign v_RM_11541_out0 = v_RM_3470_out0;
assign v_RM_11543_out0 = v_RM_3471_out0;
assign v_RM_11545_out0 = v_RM_3472_out0;
assign v_RM_11547_out0 = v_RM_3473_out0;
assign v_RM_11982_out0 = v_RM_3683_out0;
assign v_RM_11984_out0 = v_RM_3684_out0;
assign v_RM_11988_out0 = v_RM_3686_out0;
assign v_RM_11990_out0 = v_RM_3687_out0;
assign v_RM_11992_out0 = v_RM_3688_out0;
assign v_RM_11995_out0 = v_RM_3689_out0;
assign v_RM_11997_out0 = v_RM_3690_out0;
assign v_RM_11999_out0 = v_RM_3691_out0;
assign v_RM_12001_out0 = v_RM_3692_out0;
assign v_RM_12003_out0 = v_RM_3693_out0;
assign v_RM_12005_out0 = v_RM_3694_out0;
assign v_RM_12007_out0 = v_RM_3695_out0;
assign v_RM_12009_out0 = v_RM_3696_out0;
assign v_RM_12011_out0 = v_RM_3697_out0;
assign v_G2_12481_out0 = v_RD_6090_out0 && v_RM_11530_out0;
assign v_G2_12945_out0 = v_RD_6554_out0 && v_RM_11994_out0;
assign v_CARRY_5090_out0 = v_G2_12481_out0;
assign v_CARRY_5554_out0 = v_G2_12945_out0;
assign v_G1_7933_out0 = ((v_RD_6078_out0 && !v_RM_11518_out0) || (!v_RD_6078_out0) && v_RM_11518_out0);
assign v_G1_7935_out0 = ((v_RD_6080_out0 && !v_RM_11520_out0) || (!v_RD_6080_out0) && v_RM_11520_out0);
assign v_G1_7939_out0 = ((v_RD_6084_out0 && !v_RM_11524_out0) || (!v_RD_6084_out0) && v_RM_11524_out0);
assign v_G1_7941_out0 = ((v_RD_6086_out0 && !v_RM_11526_out0) || (!v_RD_6086_out0) && v_RM_11526_out0);
assign v_G1_7943_out0 = ((v_RD_6088_out0 && !v_RM_11528_out0) || (!v_RD_6088_out0) && v_RM_11528_out0);
assign v_G1_7946_out0 = ((v_RD_6091_out0 && !v_RM_11531_out0) || (!v_RD_6091_out0) && v_RM_11531_out0);
assign v_G1_7948_out0 = ((v_RD_6093_out0 && !v_RM_11533_out0) || (!v_RD_6093_out0) && v_RM_11533_out0);
assign v_G1_7950_out0 = ((v_RD_6095_out0 && !v_RM_11535_out0) || (!v_RD_6095_out0) && v_RM_11535_out0);
assign v_G1_7952_out0 = ((v_RD_6097_out0 && !v_RM_11537_out0) || (!v_RD_6097_out0) && v_RM_11537_out0);
assign v_G1_7954_out0 = ((v_RD_6099_out0 && !v_RM_11539_out0) || (!v_RD_6099_out0) && v_RM_11539_out0);
assign v_G1_7956_out0 = ((v_RD_6101_out0 && !v_RM_11541_out0) || (!v_RD_6101_out0) && v_RM_11541_out0);
assign v_G1_7958_out0 = ((v_RD_6103_out0 && !v_RM_11543_out0) || (!v_RD_6103_out0) && v_RM_11543_out0);
assign v_G1_7960_out0 = ((v_RD_6105_out0 && !v_RM_11545_out0) || (!v_RD_6105_out0) && v_RM_11545_out0);
assign v_G1_7962_out0 = ((v_RD_6107_out0 && !v_RM_11547_out0) || (!v_RD_6107_out0) && v_RM_11547_out0);
assign v_G1_8397_out0 = ((v_RD_6542_out0 && !v_RM_11982_out0) || (!v_RD_6542_out0) && v_RM_11982_out0);
assign v_G1_8399_out0 = ((v_RD_6544_out0 && !v_RM_11984_out0) || (!v_RD_6544_out0) && v_RM_11984_out0);
assign v_G1_8403_out0 = ((v_RD_6548_out0 && !v_RM_11988_out0) || (!v_RD_6548_out0) && v_RM_11988_out0);
assign v_G1_8405_out0 = ((v_RD_6550_out0 && !v_RM_11990_out0) || (!v_RD_6550_out0) && v_RM_11990_out0);
assign v_G1_8407_out0 = ((v_RD_6552_out0 && !v_RM_11992_out0) || (!v_RD_6552_out0) && v_RM_11992_out0);
assign v_G1_8410_out0 = ((v_RD_6555_out0 && !v_RM_11995_out0) || (!v_RD_6555_out0) && v_RM_11995_out0);
assign v_G1_8412_out0 = ((v_RD_6557_out0 && !v_RM_11997_out0) || (!v_RD_6557_out0) && v_RM_11997_out0);
assign v_G1_8414_out0 = ((v_RD_6559_out0 && !v_RM_11999_out0) || (!v_RD_6559_out0) && v_RM_11999_out0);
assign v_G1_8416_out0 = ((v_RD_6561_out0 && !v_RM_12001_out0) || (!v_RD_6561_out0) && v_RM_12001_out0);
assign v_G1_8418_out0 = ((v_RD_6563_out0 && !v_RM_12003_out0) || (!v_RD_6563_out0) && v_RM_12003_out0);
assign v_G1_8420_out0 = ((v_RD_6565_out0 && !v_RM_12005_out0) || (!v_RD_6565_out0) && v_RM_12005_out0);
assign v_G1_8422_out0 = ((v_RD_6567_out0 && !v_RM_12007_out0) || (!v_RD_6567_out0) && v_RM_12007_out0);
assign v_G1_8424_out0 = ((v_RD_6569_out0 && !v_RM_12009_out0) || (!v_RD_6569_out0) && v_RM_12009_out0);
assign v_G1_8426_out0 = ((v_RD_6571_out0 && !v_RM_12011_out0) || (!v_RD_6571_out0) && v_RM_12011_out0);
assign v_S_9091_out0 = v_G1_7945_out0;
assign v_S_9555_out0 = v_G1_8409_out0;
assign v_G2_12469_out0 = v_RD_6078_out0 && v_RM_11518_out0;
assign v_G2_12471_out0 = v_RD_6080_out0 && v_RM_11520_out0;
assign v_G2_12475_out0 = v_RD_6084_out0 && v_RM_11524_out0;
assign v_G2_12477_out0 = v_RD_6086_out0 && v_RM_11526_out0;
assign v_G2_12479_out0 = v_RD_6088_out0 && v_RM_11528_out0;
assign v_G2_12482_out0 = v_RD_6091_out0 && v_RM_11531_out0;
assign v_G2_12484_out0 = v_RD_6093_out0 && v_RM_11533_out0;
assign v_G2_12486_out0 = v_RD_6095_out0 && v_RM_11535_out0;
assign v_G2_12488_out0 = v_RD_6097_out0 && v_RM_11537_out0;
assign v_G2_12490_out0 = v_RD_6099_out0 && v_RM_11539_out0;
assign v_G2_12492_out0 = v_RD_6101_out0 && v_RM_11541_out0;
assign v_G2_12494_out0 = v_RD_6103_out0 && v_RM_11543_out0;
assign v_G2_12496_out0 = v_RD_6105_out0 && v_RM_11545_out0;
assign v_G2_12498_out0 = v_RD_6107_out0 && v_RM_11547_out0;
assign v_G2_12933_out0 = v_RD_6542_out0 && v_RM_11982_out0;
assign v_G2_12935_out0 = v_RD_6544_out0 && v_RM_11984_out0;
assign v_G2_12939_out0 = v_RD_6548_out0 && v_RM_11988_out0;
assign v_G2_12941_out0 = v_RD_6550_out0 && v_RM_11990_out0;
assign v_G2_12943_out0 = v_RD_6552_out0 && v_RM_11992_out0;
assign v_G2_12946_out0 = v_RD_6555_out0 && v_RM_11995_out0;
assign v_G2_12948_out0 = v_RD_6557_out0 && v_RM_11997_out0;
assign v_G2_12950_out0 = v_RD_6559_out0 && v_RM_11999_out0;
assign v_G2_12952_out0 = v_RD_6561_out0 && v_RM_12001_out0;
assign v_G2_12954_out0 = v_RD_6563_out0 && v_RM_12003_out0;
assign v_G2_12956_out0 = v_RD_6565_out0 && v_RM_12005_out0;
assign v_G2_12958_out0 = v_RD_6567_out0 && v_RM_12007_out0;
assign v_G2_12960_out0 = v_RD_6569_out0 && v_RM_12009_out0;
assign v_G2_12962_out0 = v_RD_6571_out0 && v_RM_12011_out0;
assign v_S_4672_out0 = v_S_9091_out0;
assign v_S_4687_out0 = v_S_9555_out0;
assign v_CARRY_5078_out0 = v_G2_12469_out0;
assign v_CARRY_5080_out0 = v_G2_12471_out0;
assign v_CARRY_5084_out0 = v_G2_12475_out0;
assign v_CARRY_5086_out0 = v_G2_12477_out0;
assign v_CARRY_5088_out0 = v_G2_12479_out0;
assign v_CARRY_5091_out0 = v_G2_12482_out0;
assign v_CARRY_5093_out0 = v_G2_12484_out0;
assign v_CARRY_5095_out0 = v_G2_12486_out0;
assign v_CARRY_5097_out0 = v_G2_12488_out0;
assign v_CARRY_5099_out0 = v_G2_12490_out0;
assign v_CARRY_5101_out0 = v_G2_12492_out0;
assign v_CARRY_5103_out0 = v_G2_12494_out0;
assign v_CARRY_5105_out0 = v_G2_12496_out0;
assign v_CARRY_5107_out0 = v_G2_12498_out0;
assign v_CARRY_5542_out0 = v_G2_12933_out0;
assign v_CARRY_5544_out0 = v_G2_12935_out0;
assign v_CARRY_5548_out0 = v_G2_12939_out0;
assign v_CARRY_5550_out0 = v_G2_12941_out0;
assign v_CARRY_5552_out0 = v_G2_12943_out0;
assign v_CARRY_5555_out0 = v_G2_12946_out0;
assign v_CARRY_5557_out0 = v_G2_12948_out0;
assign v_CARRY_5559_out0 = v_G2_12950_out0;
assign v_CARRY_5561_out0 = v_G2_12952_out0;
assign v_CARRY_5563_out0 = v_G2_12954_out0;
assign v_CARRY_5565_out0 = v_G2_12956_out0;
assign v_CARRY_5567_out0 = v_G2_12958_out0;
assign v_CARRY_5569_out0 = v_G2_12960_out0;
assign v_CARRY_5571_out0 = v_G2_12962_out0;
assign v_S_9079_out0 = v_G1_7933_out0;
assign v_S_9081_out0 = v_G1_7935_out0;
assign v_S_9085_out0 = v_G1_7939_out0;
assign v_S_9087_out0 = v_G1_7941_out0;
assign v_S_9089_out0 = v_G1_7943_out0;
assign v_S_9092_out0 = v_G1_7946_out0;
assign v_S_9094_out0 = v_G1_7948_out0;
assign v_S_9096_out0 = v_G1_7950_out0;
assign v_S_9098_out0 = v_G1_7952_out0;
assign v_S_9100_out0 = v_G1_7954_out0;
assign v_S_9102_out0 = v_G1_7956_out0;
assign v_S_9104_out0 = v_G1_7958_out0;
assign v_S_9106_out0 = v_G1_7960_out0;
assign v_S_9108_out0 = v_G1_7962_out0;
assign v_S_9543_out0 = v_G1_8397_out0;
assign v_S_9545_out0 = v_G1_8399_out0;
assign v_S_9549_out0 = v_G1_8403_out0;
assign v_S_9551_out0 = v_G1_8405_out0;
assign v_S_9553_out0 = v_G1_8407_out0;
assign v_S_9556_out0 = v_G1_8410_out0;
assign v_S_9558_out0 = v_G1_8412_out0;
assign v_S_9560_out0 = v_G1_8414_out0;
assign v_S_9562_out0 = v_G1_8416_out0;
assign v_S_9564_out0 = v_G1_8418_out0;
assign v_S_9566_out0 = v_G1_8420_out0;
assign v_S_9568_out0 = v_G1_8422_out0;
assign v_S_9570_out0 = v_G1_8424_out0;
assign v_S_9572_out0 = v_G1_8426_out0;
assign v_CIN_9920_out0 = v_CARRY_5090_out0;
assign v_CIN_10144_out0 = v_CARRY_5554_out0;
assign v_RD_6096_out0 = v_CIN_9920_out0;
assign v_RD_6560_out0 = v_CIN_10144_out0;
assign v_RM_11519_out0 = v_S_9079_out0;
assign v_RM_11521_out0 = v_S_9081_out0;
assign v_RM_11525_out0 = v_S_9085_out0;
assign v_RM_11527_out0 = v_S_9087_out0;
assign v_RM_11529_out0 = v_S_9089_out0;
assign v_RM_11532_out0 = v_S_9092_out0;
assign v_RM_11534_out0 = v_S_9094_out0;
assign v_RM_11536_out0 = v_S_9096_out0;
assign v_RM_11538_out0 = v_S_9098_out0;
assign v_RM_11540_out0 = v_S_9100_out0;
assign v_RM_11542_out0 = v_S_9102_out0;
assign v_RM_11544_out0 = v_S_9104_out0;
assign v_RM_11546_out0 = v_S_9106_out0;
assign v_RM_11548_out0 = v_S_9108_out0;
assign v_RM_11983_out0 = v_S_9543_out0;
assign v_RM_11985_out0 = v_S_9545_out0;
assign v_RM_11989_out0 = v_S_9549_out0;
assign v_RM_11991_out0 = v_S_9551_out0;
assign v_RM_11993_out0 = v_S_9553_out0;
assign v_RM_11996_out0 = v_S_9556_out0;
assign v_RM_11998_out0 = v_S_9558_out0;
assign v_RM_12000_out0 = v_S_9560_out0;
assign v_RM_12002_out0 = v_S_9562_out0;
assign v_RM_12004_out0 = v_S_9564_out0;
assign v_RM_12006_out0 = v_S_9566_out0;
assign v_RM_12008_out0 = v_S_9568_out0;
assign v_RM_12010_out0 = v_S_9570_out0;
assign v_RM_12012_out0 = v_S_9572_out0;
assign v__13709_out0 = { v__10767_out0,v_S_4672_out0 };
assign v__13710_out0 = { v__10768_out0,v_S_4687_out0 };
assign v_G1_7951_out0 = ((v_RD_6096_out0 && !v_RM_11536_out0) || (!v_RD_6096_out0) && v_RM_11536_out0);
assign v_G1_8415_out0 = ((v_RD_6560_out0 && !v_RM_12000_out0) || (!v_RD_6560_out0) && v_RM_12000_out0);
assign v_G2_12487_out0 = v_RD_6096_out0 && v_RM_11536_out0;
assign v_G2_12951_out0 = v_RD_6560_out0 && v_RM_12000_out0;
assign v_CARRY_5096_out0 = v_G2_12487_out0;
assign v_CARRY_5560_out0 = v_G2_12951_out0;
assign v_S_9097_out0 = v_G1_7951_out0;
assign v_S_9561_out0 = v_G1_8415_out0;
assign v_S_1331_out0 = v_S_9097_out0;
assign v_S_1555_out0 = v_S_9561_out0;
assign v_G1_4107_out0 = v_CARRY_5096_out0 || v_CARRY_5095_out0;
assign v_G1_4331_out0 = v_CARRY_5560_out0 || v_CARRY_5559_out0;
assign v_COUT_799_out0 = v_G1_4107_out0;
assign v_COUT_1023_out0 = v_G1_4331_out0;
assign v_CIN_9926_out0 = v_COUT_799_out0;
assign v_CIN_10150_out0 = v_COUT_1023_out0;
assign v_RD_6108_out0 = v_CIN_9926_out0;
assign v_RD_6572_out0 = v_CIN_10150_out0;
assign v_G1_7963_out0 = ((v_RD_6108_out0 && !v_RM_11548_out0) || (!v_RD_6108_out0) && v_RM_11548_out0);
assign v_G1_8427_out0 = ((v_RD_6572_out0 && !v_RM_12012_out0) || (!v_RD_6572_out0) && v_RM_12012_out0);
assign v_G2_12499_out0 = v_RD_6108_out0 && v_RM_11548_out0;
assign v_G2_12963_out0 = v_RD_6572_out0 && v_RM_12012_out0;
assign v_CARRY_5108_out0 = v_G2_12499_out0;
assign v_CARRY_5572_out0 = v_G2_12963_out0;
assign v_S_9109_out0 = v_G1_7963_out0;
assign v_S_9573_out0 = v_G1_8427_out0;
assign v_S_1337_out0 = v_S_9109_out0;
assign v_S_1561_out0 = v_S_9573_out0;
assign v_G1_4113_out0 = v_CARRY_5108_out0 || v_CARRY_5107_out0;
assign v_G1_4337_out0 = v_CARRY_5572_out0 || v_CARRY_5571_out0;
assign v_COUT_805_out0 = v_G1_4113_out0;
assign v_COUT_1029_out0 = v_G1_4337_out0;
assign v__4789_out0 = { v_S_1331_out0,v_S_1337_out0 };
assign v__4804_out0 = { v_S_1555_out0,v_S_1561_out0 };
assign v_CIN_9921_out0 = v_COUT_805_out0;
assign v_CIN_10145_out0 = v_COUT_1029_out0;
assign v_RD_6098_out0 = v_CIN_9921_out0;
assign v_RD_6562_out0 = v_CIN_10145_out0;
assign v_G1_7953_out0 = ((v_RD_6098_out0 && !v_RM_11538_out0) || (!v_RD_6098_out0) && v_RM_11538_out0);
assign v_G1_8417_out0 = ((v_RD_6562_out0 && !v_RM_12002_out0) || (!v_RD_6562_out0) && v_RM_12002_out0);
assign v_G2_12489_out0 = v_RD_6098_out0 && v_RM_11538_out0;
assign v_G2_12953_out0 = v_RD_6562_out0 && v_RM_12002_out0;
assign v_CARRY_5098_out0 = v_G2_12489_out0;
assign v_CARRY_5562_out0 = v_G2_12953_out0;
assign v_S_9099_out0 = v_G1_7953_out0;
assign v_S_9563_out0 = v_G1_8417_out0;
assign v_S_1332_out0 = v_S_9099_out0;
assign v_S_1556_out0 = v_S_9563_out0;
assign v_G1_4108_out0 = v_CARRY_5098_out0 || v_CARRY_5097_out0;
assign v_G1_4332_out0 = v_CARRY_5562_out0 || v_CARRY_5561_out0;
assign v_COUT_800_out0 = v_G1_4108_out0;
assign v_COUT_1024_out0 = v_G1_4332_out0;
assign v__2559_out0 = { v__4789_out0,v_S_1332_out0 };
assign v__2574_out0 = { v__4804_out0,v_S_1556_out0 };
assign v_CIN_9916_out0 = v_COUT_800_out0;
assign v_CIN_10140_out0 = v_COUT_1024_out0;
assign v_RD_6087_out0 = v_CIN_9916_out0;
assign v_RD_6551_out0 = v_CIN_10140_out0;
assign v_G1_7942_out0 = ((v_RD_6087_out0 && !v_RM_11527_out0) || (!v_RD_6087_out0) && v_RM_11527_out0);
assign v_G1_8406_out0 = ((v_RD_6551_out0 && !v_RM_11991_out0) || (!v_RD_6551_out0) && v_RM_11991_out0);
assign v_G2_12478_out0 = v_RD_6087_out0 && v_RM_11527_out0;
assign v_G2_12942_out0 = v_RD_6551_out0 && v_RM_11991_out0;
assign v_CARRY_5087_out0 = v_G2_12478_out0;
assign v_CARRY_5551_out0 = v_G2_12942_out0;
assign v_S_9088_out0 = v_G1_7942_out0;
assign v_S_9552_out0 = v_G1_8406_out0;
assign v_S_1327_out0 = v_S_9088_out0;
assign v_S_1551_out0 = v_S_9552_out0;
assign v_G1_4103_out0 = v_CARRY_5087_out0 || v_CARRY_5086_out0;
assign v_G1_4327_out0 = v_CARRY_5551_out0 || v_CARRY_5550_out0;
assign v_COUT_795_out0 = v_G1_4103_out0;
assign v_COUT_1019_out0 = v_G1_4327_out0;
assign v__7039_out0 = { v__2559_out0,v_S_1327_out0 };
assign v__7054_out0 = { v__2574_out0,v_S_1551_out0 };
assign v_CIN_9915_out0 = v_COUT_795_out0;
assign v_CIN_10139_out0 = v_COUT_1019_out0;
assign v_RD_6085_out0 = v_CIN_9915_out0;
assign v_RD_6549_out0 = v_CIN_10139_out0;
assign v_G1_7940_out0 = ((v_RD_6085_out0 && !v_RM_11525_out0) || (!v_RD_6085_out0) && v_RM_11525_out0);
assign v_G1_8404_out0 = ((v_RD_6549_out0 && !v_RM_11989_out0) || (!v_RD_6549_out0) && v_RM_11989_out0);
assign v_G2_12476_out0 = v_RD_6085_out0 && v_RM_11525_out0;
assign v_G2_12940_out0 = v_RD_6549_out0 && v_RM_11989_out0;
assign v_CARRY_5085_out0 = v_G2_12476_out0;
assign v_CARRY_5549_out0 = v_G2_12940_out0;
assign v_S_9086_out0 = v_G1_7940_out0;
assign v_S_9550_out0 = v_G1_8404_out0;
assign v_S_1326_out0 = v_S_9086_out0;
assign v_S_1550_out0 = v_S_9550_out0;
assign v_G1_4102_out0 = v_CARRY_5085_out0 || v_CARRY_5084_out0;
assign v_G1_4326_out0 = v_CARRY_5549_out0 || v_CARRY_5548_out0;
assign v_COUT_794_out0 = v_G1_4102_out0;
assign v_COUT_1018_out0 = v_G1_4326_out0;
assign v__13525_out0 = { v__7039_out0,v_S_1326_out0 };
assign v__13540_out0 = { v__7054_out0,v_S_1550_out0 };
assign v_CIN_9922_out0 = v_COUT_794_out0;
assign v_CIN_10146_out0 = v_COUT_1018_out0;
assign v_RD_6100_out0 = v_CIN_9922_out0;
assign v_RD_6564_out0 = v_CIN_10146_out0;
assign v_G1_7955_out0 = ((v_RD_6100_out0 && !v_RM_11540_out0) || (!v_RD_6100_out0) && v_RM_11540_out0);
assign v_G1_8419_out0 = ((v_RD_6564_out0 && !v_RM_12004_out0) || (!v_RD_6564_out0) && v_RM_12004_out0);
assign v_G2_12491_out0 = v_RD_6100_out0 && v_RM_11540_out0;
assign v_G2_12955_out0 = v_RD_6564_out0 && v_RM_12004_out0;
assign v_CARRY_5100_out0 = v_G2_12491_out0;
assign v_CARRY_5564_out0 = v_G2_12955_out0;
assign v_S_9101_out0 = v_G1_7955_out0;
assign v_S_9565_out0 = v_G1_8419_out0;
assign v_S_1333_out0 = v_S_9101_out0;
assign v_S_1557_out0 = v_S_9565_out0;
assign v_G1_4109_out0 = v_CARRY_5100_out0 || v_CARRY_5099_out0;
assign v_G1_4333_out0 = v_CARRY_5564_out0 || v_CARRY_5563_out0;
assign v_COUT_801_out0 = v_G1_4109_out0;
assign v_COUT_1025_out0 = v_G1_4333_out0;
assign v__3318_out0 = { v__13525_out0,v_S_1333_out0 };
assign v__3333_out0 = { v__13540_out0,v_S_1557_out0 };
assign v_CIN_9923_out0 = v_COUT_801_out0;
assign v_CIN_10147_out0 = v_COUT_1025_out0;
assign v_RD_6102_out0 = v_CIN_9923_out0;
assign v_RD_6566_out0 = v_CIN_10147_out0;
assign v_G1_7957_out0 = ((v_RD_6102_out0 && !v_RM_11542_out0) || (!v_RD_6102_out0) && v_RM_11542_out0);
assign v_G1_8421_out0 = ((v_RD_6566_out0 && !v_RM_12006_out0) || (!v_RD_6566_out0) && v_RM_12006_out0);
assign v_G2_12493_out0 = v_RD_6102_out0 && v_RM_11542_out0;
assign v_G2_12957_out0 = v_RD_6566_out0 && v_RM_12006_out0;
assign v_CARRY_5102_out0 = v_G2_12493_out0;
assign v_CARRY_5566_out0 = v_G2_12957_out0;
assign v_S_9103_out0 = v_G1_7957_out0;
assign v_S_9567_out0 = v_G1_8421_out0;
assign v_S_1334_out0 = v_S_9103_out0;
assign v_S_1558_out0 = v_S_9567_out0;
assign v_G1_4110_out0 = v_CARRY_5102_out0 || v_CARRY_5101_out0;
assign v_G1_4334_out0 = v_CARRY_5566_out0 || v_CARRY_5565_out0;
assign v_COUT_802_out0 = v_G1_4110_out0;
assign v_COUT_1026_out0 = v_G1_4334_out0;
assign v__7154_out0 = { v__3318_out0,v_S_1334_out0 };
assign v__7169_out0 = { v__3333_out0,v_S_1558_out0 };
assign v_CIN_9925_out0 = v_COUT_802_out0;
assign v_CIN_10149_out0 = v_COUT_1026_out0;
assign v_RD_6106_out0 = v_CIN_9925_out0;
assign v_RD_6570_out0 = v_CIN_10149_out0;
assign v_G1_7961_out0 = ((v_RD_6106_out0 && !v_RM_11546_out0) || (!v_RD_6106_out0) && v_RM_11546_out0);
assign v_G1_8425_out0 = ((v_RD_6570_out0 && !v_RM_12010_out0) || (!v_RD_6570_out0) && v_RM_12010_out0);
assign v_G2_12497_out0 = v_RD_6106_out0 && v_RM_11546_out0;
assign v_G2_12961_out0 = v_RD_6570_out0 && v_RM_12010_out0;
assign v_CARRY_5106_out0 = v_G2_12497_out0;
assign v_CARRY_5570_out0 = v_G2_12961_out0;
assign v_S_9107_out0 = v_G1_7961_out0;
assign v_S_9571_out0 = v_G1_8425_out0;
assign v_S_1336_out0 = v_S_9107_out0;
assign v_S_1560_out0 = v_S_9571_out0;
assign v_G1_4112_out0 = v_CARRY_5106_out0 || v_CARRY_5105_out0;
assign v_G1_4336_out0 = v_CARRY_5570_out0 || v_CARRY_5569_out0;
assign v_COUT_804_out0 = v_G1_4112_out0;
assign v_COUT_1028_out0 = v_G1_4336_out0;
assign v__4756_out0 = { v__7154_out0,v_S_1336_out0 };
assign v__4771_out0 = { v__7169_out0,v_S_1560_out0 };
assign v_CIN_9918_out0 = v_COUT_804_out0;
assign v_CIN_10142_out0 = v_COUT_1028_out0;
assign v_RD_6092_out0 = v_CIN_9918_out0;
assign v_RD_6556_out0 = v_CIN_10142_out0;
assign v_G1_7947_out0 = ((v_RD_6092_out0 && !v_RM_11532_out0) || (!v_RD_6092_out0) && v_RM_11532_out0);
assign v_G1_8411_out0 = ((v_RD_6556_out0 && !v_RM_11996_out0) || (!v_RD_6556_out0) && v_RM_11996_out0);
assign v_G2_12483_out0 = v_RD_6092_out0 && v_RM_11532_out0;
assign v_G2_12947_out0 = v_RD_6556_out0 && v_RM_11996_out0;
assign v_CARRY_5092_out0 = v_G2_12483_out0;
assign v_CARRY_5556_out0 = v_G2_12947_out0;
assign v_S_9093_out0 = v_G1_7947_out0;
assign v_S_9557_out0 = v_G1_8411_out0;
assign v_S_1329_out0 = v_S_9093_out0;
assign v_S_1553_out0 = v_S_9557_out0;
assign v_G1_4105_out0 = v_CARRY_5092_out0 || v_CARRY_5091_out0;
assign v_G1_4329_out0 = v_CARRY_5556_out0 || v_CARRY_5555_out0;
assign v_COUT_797_out0 = v_G1_4105_out0;
assign v_COUT_1021_out0 = v_G1_4329_out0;
assign v__6933_out0 = { v__4756_out0,v_S_1329_out0 };
assign v__6948_out0 = { v__4771_out0,v_S_1553_out0 };
assign v_CIN_9919_out0 = v_COUT_797_out0;
assign v_CIN_10143_out0 = v_COUT_1021_out0;
assign v_RD_6094_out0 = v_CIN_9919_out0;
assign v_RD_6558_out0 = v_CIN_10143_out0;
assign v_G1_7949_out0 = ((v_RD_6094_out0 && !v_RM_11534_out0) || (!v_RD_6094_out0) && v_RM_11534_out0);
assign v_G1_8413_out0 = ((v_RD_6558_out0 && !v_RM_11998_out0) || (!v_RD_6558_out0) && v_RM_11998_out0);
assign v_G2_12485_out0 = v_RD_6094_out0 && v_RM_11534_out0;
assign v_G2_12949_out0 = v_RD_6558_out0 && v_RM_11998_out0;
assign v_CARRY_5094_out0 = v_G2_12485_out0;
assign v_CARRY_5558_out0 = v_G2_12949_out0;
assign v_S_9095_out0 = v_G1_7949_out0;
assign v_S_9559_out0 = v_G1_8413_out0;
assign v_S_1330_out0 = v_S_9095_out0;
assign v_S_1554_out0 = v_S_9559_out0;
assign v_G1_4106_out0 = v_CARRY_5094_out0 || v_CARRY_5093_out0;
assign v_G1_4330_out0 = v_CARRY_5558_out0 || v_CARRY_5557_out0;
assign v_COUT_798_out0 = v_G1_4106_out0;
assign v_COUT_1022_out0 = v_G1_4330_out0;
assign v__5809_out0 = { v__6933_out0,v_S_1330_out0 };
assign v__5824_out0 = { v__6948_out0,v_S_1554_out0 };
assign v_CIN_9924_out0 = v_COUT_798_out0;
assign v_CIN_10148_out0 = v_COUT_1022_out0;
assign v_RD_6104_out0 = v_CIN_9924_out0;
assign v_RD_6568_out0 = v_CIN_10148_out0;
assign v_G1_7959_out0 = ((v_RD_6104_out0 && !v_RM_11544_out0) || (!v_RD_6104_out0) && v_RM_11544_out0);
assign v_G1_8423_out0 = ((v_RD_6568_out0 && !v_RM_12008_out0) || (!v_RD_6568_out0) && v_RM_12008_out0);
assign v_G2_12495_out0 = v_RD_6104_out0 && v_RM_11544_out0;
assign v_G2_12959_out0 = v_RD_6568_out0 && v_RM_12008_out0;
assign v_CARRY_5104_out0 = v_G2_12495_out0;
assign v_CARRY_5568_out0 = v_G2_12959_out0;
assign v_S_9105_out0 = v_G1_7959_out0;
assign v_S_9569_out0 = v_G1_8423_out0;
assign v_S_1335_out0 = v_S_9105_out0;
assign v_S_1559_out0 = v_S_9569_out0;
assign v_G1_4111_out0 = v_CARRY_5104_out0 || v_CARRY_5103_out0;
assign v_G1_4335_out0 = v_CARRY_5568_out0 || v_CARRY_5567_out0;
assign v_COUT_803_out0 = v_G1_4111_out0;
assign v_COUT_1027_out0 = v_G1_4335_out0;
assign v__2033_out0 = { v__5809_out0,v_S_1335_out0 };
assign v__2048_out0 = { v__5824_out0,v_S_1559_out0 };
assign v_CIN_9912_out0 = v_COUT_803_out0;
assign v_CIN_10136_out0 = v_COUT_1027_out0;
assign v_RD_6079_out0 = v_CIN_9912_out0;
assign v_RD_6543_out0 = v_CIN_10136_out0;
assign v_G1_7934_out0 = ((v_RD_6079_out0 && !v_RM_11519_out0) || (!v_RD_6079_out0) && v_RM_11519_out0);
assign v_G1_8398_out0 = ((v_RD_6543_out0 && !v_RM_11983_out0) || (!v_RD_6543_out0) && v_RM_11983_out0);
assign v_G2_12470_out0 = v_RD_6079_out0 && v_RM_11519_out0;
assign v_G2_12934_out0 = v_RD_6543_out0 && v_RM_11983_out0;
assign v_CARRY_5079_out0 = v_G2_12470_out0;
assign v_CARRY_5543_out0 = v_G2_12934_out0;
assign v_S_9080_out0 = v_G1_7934_out0;
assign v_S_9544_out0 = v_G1_8398_out0;
assign v_S_1323_out0 = v_S_9080_out0;
assign v_S_1547_out0 = v_S_9544_out0;
assign v_G1_4099_out0 = v_CARRY_5079_out0 || v_CARRY_5078_out0;
assign v_G1_4323_out0 = v_CARRY_5543_out0 || v_CARRY_5542_out0;
assign v_COUT_791_out0 = v_G1_4099_out0;
assign v_COUT_1015_out0 = v_G1_4323_out0;
assign v__2800_out0 = { v__2033_out0,v_S_1323_out0 };
assign v__2815_out0 = { v__2048_out0,v_S_1547_out0 };
assign v_CIN_9917_out0 = v_COUT_791_out0;
assign v_CIN_10141_out0 = v_COUT_1015_out0;
assign v_RD_6089_out0 = v_CIN_9917_out0;
assign v_RD_6553_out0 = v_CIN_10141_out0;
assign v_G1_7944_out0 = ((v_RD_6089_out0 && !v_RM_11529_out0) || (!v_RD_6089_out0) && v_RM_11529_out0);
assign v_G1_8408_out0 = ((v_RD_6553_out0 && !v_RM_11993_out0) || (!v_RD_6553_out0) && v_RM_11993_out0);
assign v_G2_12480_out0 = v_RD_6089_out0 && v_RM_11529_out0;
assign v_G2_12944_out0 = v_RD_6553_out0 && v_RM_11993_out0;
assign v_CARRY_5089_out0 = v_G2_12480_out0;
assign v_CARRY_5553_out0 = v_G2_12944_out0;
assign v_S_9090_out0 = v_G1_7944_out0;
assign v_S_9554_out0 = v_G1_8408_out0;
assign v_S_1328_out0 = v_S_9090_out0;
assign v_S_1552_out0 = v_S_9554_out0;
assign v_G1_4104_out0 = v_CARRY_5089_out0 || v_CARRY_5088_out0;
assign v_G1_4328_out0 = v_CARRY_5553_out0 || v_CARRY_5552_out0;
assign v_COUT_796_out0 = v_G1_4104_out0;
assign v_COUT_1020_out0 = v_G1_4328_out0;
assign v__1832_out0 = { v__2800_out0,v_S_1328_out0 };
assign v__1847_out0 = { v__2815_out0,v_S_1552_out0 };
assign v_CIN_9913_out0 = v_COUT_796_out0;
assign v_CIN_10137_out0 = v_COUT_1020_out0;
assign v_RD_6081_out0 = v_CIN_9913_out0;
assign v_RD_6545_out0 = v_CIN_10137_out0;
assign v_G1_7936_out0 = ((v_RD_6081_out0 && !v_RM_11521_out0) || (!v_RD_6081_out0) && v_RM_11521_out0);
assign v_G1_8400_out0 = ((v_RD_6545_out0 && !v_RM_11985_out0) || (!v_RD_6545_out0) && v_RM_11985_out0);
assign v_G2_12472_out0 = v_RD_6081_out0 && v_RM_11521_out0;
assign v_G2_12936_out0 = v_RD_6545_out0 && v_RM_11985_out0;
assign v_CARRY_5081_out0 = v_G2_12472_out0;
assign v_CARRY_5545_out0 = v_G2_12936_out0;
assign v_S_9082_out0 = v_G1_7936_out0;
assign v_S_9546_out0 = v_G1_8400_out0;
assign v_S_1324_out0 = v_S_9082_out0;
assign v_S_1548_out0 = v_S_9546_out0;
assign v_G1_4100_out0 = v_CARRY_5081_out0 || v_CARRY_5080_out0;
assign v_G1_4324_out0 = v_CARRY_5545_out0 || v_CARRY_5544_out0;
assign v_COUT_792_out0 = v_G1_4100_out0;
assign v_COUT_1016_out0 = v_G1_4324_out0;
assign v__4556_out0 = { v__1832_out0,v_S_1324_out0 };
assign v__4571_out0 = { v__1847_out0,v_S_1548_out0 };
assign v_RM_3461_out0 = v_COUT_792_out0;
assign v_RM_3685_out0 = v_COUT_1016_out0;
assign v_RM_11522_out0 = v_RM_3461_out0;
assign v_RM_11986_out0 = v_RM_3685_out0;
assign v_G1_7937_out0 = ((v_RD_6082_out0 && !v_RM_11522_out0) || (!v_RD_6082_out0) && v_RM_11522_out0);
assign v_G1_8401_out0 = ((v_RD_6546_out0 && !v_RM_11986_out0) || (!v_RD_6546_out0) && v_RM_11986_out0);
assign v_G2_12473_out0 = v_RD_6082_out0 && v_RM_11522_out0;
assign v_G2_12937_out0 = v_RD_6546_out0 && v_RM_11986_out0;
assign v_CARRY_5082_out0 = v_G2_12473_out0;
assign v_CARRY_5546_out0 = v_G2_12937_out0;
assign v_S_9083_out0 = v_G1_7937_out0;
assign v_S_9547_out0 = v_G1_8401_out0;
assign v_RM_11523_out0 = v_S_9083_out0;
assign v_RM_11987_out0 = v_S_9547_out0;
assign v_G1_7938_out0 = ((v_RD_6083_out0 && !v_RM_11523_out0) || (!v_RD_6083_out0) && v_RM_11523_out0);
assign v_G1_8402_out0 = ((v_RD_6547_out0 && !v_RM_11987_out0) || (!v_RD_6547_out0) && v_RM_11987_out0);
assign v_G2_12474_out0 = v_RD_6083_out0 && v_RM_11523_out0;
assign v_G2_12938_out0 = v_RD_6547_out0 && v_RM_11987_out0;
assign v_CARRY_5083_out0 = v_G2_12474_out0;
assign v_CARRY_5547_out0 = v_G2_12938_out0;
assign v_S_9084_out0 = v_G1_7938_out0;
assign v_S_9548_out0 = v_G1_8402_out0;
assign v_S_1325_out0 = v_S_9084_out0;
assign v_S_1549_out0 = v_S_9548_out0;
assign v_G1_4101_out0 = v_CARRY_5083_out0 || v_CARRY_5082_out0;
assign v_G1_4325_out0 = v_CARRY_5547_out0 || v_CARRY_5546_out0;
assign v_COUT_793_out0 = v_G1_4101_out0;
assign v_COUT_1017_out0 = v_G1_4325_out0;
assign v__10658_out0 = { v__4556_out0,v_S_1325_out0 };
assign v__10673_out0 = { v__4571_out0,v_S_1549_out0 };
assign v__10953_out0 = { v__10658_out0,v_COUT_793_out0 };
assign v__10968_out0 = { v__10673_out0,v_COUT_1017_out0 };
assign v_COUT_10923_out0 = v__10953_out0;
assign v_COUT_10938_out0 = v__10968_out0;
assign v_CIN_2361_out0 = v_COUT_10923_out0;
assign v_CIN_2376_out0 = v_COUT_10938_out0;
assign v__474_out0 = v_CIN_2361_out0[8:8];
assign v__489_out0 = v_CIN_2376_out0[8:8];
assign v__1779_out0 = v_CIN_2361_out0[6:6];
assign v__1794_out0 = v_CIN_2376_out0[6:6];
assign v__2161_out0 = v_CIN_2361_out0[3:3];
assign v__2176_out0 = v_CIN_2376_out0[3:3];
assign v__2200_out0 = v_CIN_2361_out0[15:15];
assign v__2214_out0 = v_CIN_2376_out0[15:15];
assign v__2508_out0 = v_CIN_2361_out0[0:0];
assign v__2523_out0 = v_CIN_2376_out0[0:0];
assign v__3057_out0 = v_CIN_2361_out0[9:9];
assign v__3072_out0 = v_CIN_2376_out0[9:9];
assign v__3091_out0 = v_CIN_2361_out0[2:2];
assign v__3106_out0 = v_CIN_2376_out0[2:2];
assign v__3145_out0 = v_CIN_2361_out0[7:7];
assign v__3160_out0 = v_CIN_2376_out0[7:7];
assign v__3829_out0 = v_CIN_2361_out0[1:1];
assign v__3844_out0 = v_CIN_2376_out0[1:1];
assign v__3867_out0 = v_CIN_2361_out0[10:10];
assign v__3882_out0 = v_CIN_2376_out0[10:10];
assign v__6806_out0 = v_CIN_2361_out0[11:11];
assign v__6821_out0 = v_CIN_2376_out0[11:11];
assign v__7650_out0 = v_CIN_2361_out0[12:12];
assign v__7665_out0 = v_CIN_2376_out0[12:12];
assign v__8705_out0 = v_CIN_2361_out0[13:13];
assign v__8720_out0 = v_CIN_2376_out0[13:13];
assign v__8775_out0 = v_CIN_2361_out0[14:14];
assign v__8790_out0 = v_CIN_2376_out0[14:14];
assign v__10725_out0 = v_CIN_2361_out0[5:5];
assign v__10740_out0 = v_CIN_2376_out0[5:5];
assign v__13454_out0 = v_CIN_2361_out0[4:4];
assign v__13469_out0 = v_CIN_2376_out0[4:4];
assign v_RM_3444_out0 = v__7650_out0;
assign v_RM_3445_out0 = v__8775_out0;
assign v_RM_3447_out0 = v__10725_out0;
assign v_RM_3448_out0 = v__13454_out0;
assign v_RM_3449_out0 = v__8705_out0;
assign v_RM_3450_out0 = v__3057_out0;
assign v_RM_3451_out0 = v__3867_out0;
assign v_RM_3452_out0 = v__3829_out0;
assign v_RM_3453_out0 = v__2161_out0;
assign v_RM_3454_out0 = v__1779_out0;
assign v_RM_3455_out0 = v__3145_out0;
assign v_RM_3456_out0 = v__6806_out0;
assign v_RM_3457_out0 = v__474_out0;
assign v_RM_3458_out0 = v__3091_out0;
assign v_RM_3668_out0 = v__7665_out0;
assign v_RM_3669_out0 = v__8790_out0;
assign v_RM_3671_out0 = v__10740_out0;
assign v_RM_3672_out0 = v__13469_out0;
assign v_RM_3673_out0 = v__8720_out0;
assign v_RM_3674_out0 = v__3072_out0;
assign v_RM_3675_out0 = v__3882_out0;
assign v_RM_3676_out0 = v__3844_out0;
assign v_RM_3677_out0 = v__2176_out0;
assign v_RM_3678_out0 = v__1794_out0;
assign v_RM_3679_out0 = v__3160_out0;
assign v_RM_3680_out0 = v__6821_out0;
assign v_RM_3681_out0 = v__489_out0;
assign v_RM_3682_out0 = v__3106_out0;
assign v_CIN_9899_out0 = v__2200_out0;
assign v_CIN_10123_out0 = v__2214_out0;
assign v_RM_11499_out0 = v__2508_out0;
assign v_RM_11963_out0 = v__2523_out0;
assign v_RD_6052_out0 = v_CIN_9899_out0;
assign v_RD_6516_out0 = v_CIN_10123_out0;
assign v_G1_7914_out0 = ((v_RD_6059_out0 && !v_RM_11499_out0) || (!v_RD_6059_out0) && v_RM_11499_out0);
assign v_G1_8378_out0 = ((v_RD_6523_out0 && !v_RM_11963_out0) || (!v_RD_6523_out0) && v_RM_11963_out0);
assign v_RM_11487_out0 = v_RM_3444_out0;
assign v_RM_11489_out0 = v_RM_3445_out0;
assign v_RM_11493_out0 = v_RM_3447_out0;
assign v_RM_11495_out0 = v_RM_3448_out0;
assign v_RM_11497_out0 = v_RM_3449_out0;
assign v_RM_11500_out0 = v_RM_3450_out0;
assign v_RM_11502_out0 = v_RM_3451_out0;
assign v_RM_11504_out0 = v_RM_3452_out0;
assign v_RM_11506_out0 = v_RM_3453_out0;
assign v_RM_11508_out0 = v_RM_3454_out0;
assign v_RM_11510_out0 = v_RM_3455_out0;
assign v_RM_11512_out0 = v_RM_3456_out0;
assign v_RM_11514_out0 = v_RM_3457_out0;
assign v_RM_11516_out0 = v_RM_3458_out0;
assign v_RM_11951_out0 = v_RM_3668_out0;
assign v_RM_11953_out0 = v_RM_3669_out0;
assign v_RM_11957_out0 = v_RM_3671_out0;
assign v_RM_11959_out0 = v_RM_3672_out0;
assign v_RM_11961_out0 = v_RM_3673_out0;
assign v_RM_11964_out0 = v_RM_3674_out0;
assign v_RM_11966_out0 = v_RM_3675_out0;
assign v_RM_11968_out0 = v_RM_3676_out0;
assign v_RM_11970_out0 = v_RM_3677_out0;
assign v_RM_11972_out0 = v_RM_3678_out0;
assign v_RM_11974_out0 = v_RM_3679_out0;
assign v_RM_11976_out0 = v_RM_3680_out0;
assign v_RM_11978_out0 = v_RM_3681_out0;
assign v_RM_11980_out0 = v_RM_3682_out0;
assign v_G2_12450_out0 = v_RD_6059_out0 && v_RM_11499_out0;
assign v_G2_12914_out0 = v_RD_6523_out0 && v_RM_11963_out0;
assign v_CARRY_5059_out0 = v_G2_12450_out0;
assign v_CARRY_5523_out0 = v_G2_12914_out0;
assign v_G1_7902_out0 = ((v_RD_6047_out0 && !v_RM_11487_out0) || (!v_RD_6047_out0) && v_RM_11487_out0);
assign v_G1_7904_out0 = ((v_RD_6049_out0 && !v_RM_11489_out0) || (!v_RD_6049_out0) && v_RM_11489_out0);
assign v_G1_7908_out0 = ((v_RD_6053_out0 && !v_RM_11493_out0) || (!v_RD_6053_out0) && v_RM_11493_out0);
assign v_G1_7910_out0 = ((v_RD_6055_out0 && !v_RM_11495_out0) || (!v_RD_6055_out0) && v_RM_11495_out0);
assign v_G1_7912_out0 = ((v_RD_6057_out0 && !v_RM_11497_out0) || (!v_RD_6057_out0) && v_RM_11497_out0);
assign v_G1_7915_out0 = ((v_RD_6060_out0 && !v_RM_11500_out0) || (!v_RD_6060_out0) && v_RM_11500_out0);
assign v_G1_7917_out0 = ((v_RD_6062_out0 && !v_RM_11502_out0) || (!v_RD_6062_out0) && v_RM_11502_out0);
assign v_G1_7919_out0 = ((v_RD_6064_out0 && !v_RM_11504_out0) || (!v_RD_6064_out0) && v_RM_11504_out0);
assign v_G1_7921_out0 = ((v_RD_6066_out0 && !v_RM_11506_out0) || (!v_RD_6066_out0) && v_RM_11506_out0);
assign v_G1_7923_out0 = ((v_RD_6068_out0 && !v_RM_11508_out0) || (!v_RD_6068_out0) && v_RM_11508_out0);
assign v_G1_7925_out0 = ((v_RD_6070_out0 && !v_RM_11510_out0) || (!v_RD_6070_out0) && v_RM_11510_out0);
assign v_G1_7927_out0 = ((v_RD_6072_out0 && !v_RM_11512_out0) || (!v_RD_6072_out0) && v_RM_11512_out0);
assign v_G1_7929_out0 = ((v_RD_6074_out0 && !v_RM_11514_out0) || (!v_RD_6074_out0) && v_RM_11514_out0);
assign v_G1_7931_out0 = ((v_RD_6076_out0 && !v_RM_11516_out0) || (!v_RD_6076_out0) && v_RM_11516_out0);
assign v_G1_8366_out0 = ((v_RD_6511_out0 && !v_RM_11951_out0) || (!v_RD_6511_out0) && v_RM_11951_out0);
assign v_G1_8368_out0 = ((v_RD_6513_out0 && !v_RM_11953_out0) || (!v_RD_6513_out0) && v_RM_11953_out0);
assign v_G1_8372_out0 = ((v_RD_6517_out0 && !v_RM_11957_out0) || (!v_RD_6517_out0) && v_RM_11957_out0);
assign v_G1_8374_out0 = ((v_RD_6519_out0 && !v_RM_11959_out0) || (!v_RD_6519_out0) && v_RM_11959_out0);
assign v_G1_8376_out0 = ((v_RD_6521_out0 && !v_RM_11961_out0) || (!v_RD_6521_out0) && v_RM_11961_out0);
assign v_G1_8379_out0 = ((v_RD_6524_out0 && !v_RM_11964_out0) || (!v_RD_6524_out0) && v_RM_11964_out0);
assign v_G1_8381_out0 = ((v_RD_6526_out0 && !v_RM_11966_out0) || (!v_RD_6526_out0) && v_RM_11966_out0);
assign v_G1_8383_out0 = ((v_RD_6528_out0 && !v_RM_11968_out0) || (!v_RD_6528_out0) && v_RM_11968_out0);
assign v_G1_8385_out0 = ((v_RD_6530_out0 && !v_RM_11970_out0) || (!v_RD_6530_out0) && v_RM_11970_out0);
assign v_G1_8387_out0 = ((v_RD_6532_out0 && !v_RM_11972_out0) || (!v_RD_6532_out0) && v_RM_11972_out0);
assign v_G1_8389_out0 = ((v_RD_6534_out0 && !v_RM_11974_out0) || (!v_RD_6534_out0) && v_RM_11974_out0);
assign v_G1_8391_out0 = ((v_RD_6536_out0 && !v_RM_11976_out0) || (!v_RD_6536_out0) && v_RM_11976_out0);
assign v_G1_8393_out0 = ((v_RD_6538_out0 && !v_RM_11978_out0) || (!v_RD_6538_out0) && v_RM_11978_out0);
assign v_G1_8395_out0 = ((v_RD_6540_out0 && !v_RM_11980_out0) || (!v_RD_6540_out0) && v_RM_11980_out0);
assign v_S_9060_out0 = v_G1_7914_out0;
assign v_S_9524_out0 = v_G1_8378_out0;
assign v_G2_12438_out0 = v_RD_6047_out0 && v_RM_11487_out0;
assign v_G2_12440_out0 = v_RD_6049_out0 && v_RM_11489_out0;
assign v_G2_12444_out0 = v_RD_6053_out0 && v_RM_11493_out0;
assign v_G2_12446_out0 = v_RD_6055_out0 && v_RM_11495_out0;
assign v_G2_12448_out0 = v_RD_6057_out0 && v_RM_11497_out0;
assign v_G2_12451_out0 = v_RD_6060_out0 && v_RM_11500_out0;
assign v_G2_12453_out0 = v_RD_6062_out0 && v_RM_11502_out0;
assign v_G2_12455_out0 = v_RD_6064_out0 && v_RM_11504_out0;
assign v_G2_12457_out0 = v_RD_6066_out0 && v_RM_11506_out0;
assign v_G2_12459_out0 = v_RD_6068_out0 && v_RM_11508_out0;
assign v_G2_12461_out0 = v_RD_6070_out0 && v_RM_11510_out0;
assign v_G2_12463_out0 = v_RD_6072_out0 && v_RM_11512_out0;
assign v_G2_12465_out0 = v_RD_6074_out0 && v_RM_11514_out0;
assign v_G2_12467_out0 = v_RD_6076_out0 && v_RM_11516_out0;
assign v_G2_12902_out0 = v_RD_6511_out0 && v_RM_11951_out0;
assign v_G2_12904_out0 = v_RD_6513_out0 && v_RM_11953_out0;
assign v_G2_12908_out0 = v_RD_6517_out0 && v_RM_11957_out0;
assign v_G2_12910_out0 = v_RD_6519_out0 && v_RM_11959_out0;
assign v_G2_12912_out0 = v_RD_6521_out0 && v_RM_11961_out0;
assign v_G2_12915_out0 = v_RD_6524_out0 && v_RM_11964_out0;
assign v_G2_12917_out0 = v_RD_6526_out0 && v_RM_11966_out0;
assign v_G2_12919_out0 = v_RD_6528_out0 && v_RM_11968_out0;
assign v_G2_12921_out0 = v_RD_6530_out0 && v_RM_11970_out0;
assign v_G2_12923_out0 = v_RD_6532_out0 && v_RM_11972_out0;
assign v_G2_12925_out0 = v_RD_6534_out0 && v_RM_11974_out0;
assign v_G2_12927_out0 = v_RD_6536_out0 && v_RM_11976_out0;
assign v_G2_12929_out0 = v_RD_6538_out0 && v_RM_11978_out0;
assign v_G2_12931_out0 = v_RD_6540_out0 && v_RM_11980_out0;
assign v_S_4671_out0 = v_S_9060_out0;
assign v_S_4686_out0 = v_S_9524_out0;
assign v_CARRY_5047_out0 = v_G2_12438_out0;
assign v_CARRY_5049_out0 = v_G2_12440_out0;
assign v_CARRY_5053_out0 = v_G2_12444_out0;
assign v_CARRY_5055_out0 = v_G2_12446_out0;
assign v_CARRY_5057_out0 = v_G2_12448_out0;
assign v_CARRY_5060_out0 = v_G2_12451_out0;
assign v_CARRY_5062_out0 = v_G2_12453_out0;
assign v_CARRY_5064_out0 = v_G2_12455_out0;
assign v_CARRY_5066_out0 = v_G2_12457_out0;
assign v_CARRY_5068_out0 = v_G2_12459_out0;
assign v_CARRY_5070_out0 = v_G2_12461_out0;
assign v_CARRY_5072_out0 = v_G2_12463_out0;
assign v_CARRY_5074_out0 = v_G2_12465_out0;
assign v_CARRY_5076_out0 = v_G2_12467_out0;
assign v_CARRY_5511_out0 = v_G2_12902_out0;
assign v_CARRY_5513_out0 = v_G2_12904_out0;
assign v_CARRY_5517_out0 = v_G2_12908_out0;
assign v_CARRY_5519_out0 = v_G2_12910_out0;
assign v_CARRY_5521_out0 = v_G2_12912_out0;
assign v_CARRY_5524_out0 = v_G2_12915_out0;
assign v_CARRY_5526_out0 = v_G2_12917_out0;
assign v_CARRY_5528_out0 = v_G2_12919_out0;
assign v_CARRY_5530_out0 = v_G2_12921_out0;
assign v_CARRY_5532_out0 = v_G2_12923_out0;
assign v_CARRY_5534_out0 = v_G2_12925_out0;
assign v_CARRY_5536_out0 = v_G2_12927_out0;
assign v_CARRY_5538_out0 = v_G2_12929_out0;
assign v_CARRY_5540_out0 = v_G2_12931_out0;
assign v_S_9048_out0 = v_G1_7902_out0;
assign v_S_9050_out0 = v_G1_7904_out0;
assign v_S_9054_out0 = v_G1_7908_out0;
assign v_S_9056_out0 = v_G1_7910_out0;
assign v_S_9058_out0 = v_G1_7912_out0;
assign v_S_9061_out0 = v_G1_7915_out0;
assign v_S_9063_out0 = v_G1_7917_out0;
assign v_S_9065_out0 = v_G1_7919_out0;
assign v_S_9067_out0 = v_G1_7921_out0;
assign v_S_9069_out0 = v_G1_7923_out0;
assign v_S_9071_out0 = v_G1_7925_out0;
assign v_S_9073_out0 = v_G1_7927_out0;
assign v_S_9075_out0 = v_G1_7929_out0;
assign v_S_9077_out0 = v_G1_7931_out0;
assign v_S_9512_out0 = v_G1_8366_out0;
assign v_S_9514_out0 = v_G1_8368_out0;
assign v_S_9518_out0 = v_G1_8372_out0;
assign v_S_9520_out0 = v_G1_8374_out0;
assign v_S_9522_out0 = v_G1_8376_out0;
assign v_S_9525_out0 = v_G1_8379_out0;
assign v_S_9527_out0 = v_G1_8381_out0;
assign v_S_9529_out0 = v_G1_8383_out0;
assign v_S_9531_out0 = v_G1_8385_out0;
assign v_S_9533_out0 = v_G1_8387_out0;
assign v_S_9535_out0 = v_G1_8389_out0;
assign v_S_9537_out0 = v_G1_8391_out0;
assign v_S_9539_out0 = v_G1_8393_out0;
assign v_S_9541_out0 = v_G1_8395_out0;
assign v_CIN_9905_out0 = v_CARRY_5059_out0;
assign v_CIN_10129_out0 = v_CARRY_5523_out0;
assign v__403_out0 = { v__13709_out0,v_S_4671_out0 };
assign v__404_out0 = { v__13710_out0,v_S_4686_out0 };
assign v_RD_6065_out0 = v_CIN_9905_out0;
assign v_RD_6529_out0 = v_CIN_10129_out0;
assign v_RM_11488_out0 = v_S_9048_out0;
assign v_RM_11490_out0 = v_S_9050_out0;
assign v_RM_11494_out0 = v_S_9054_out0;
assign v_RM_11496_out0 = v_S_9056_out0;
assign v_RM_11498_out0 = v_S_9058_out0;
assign v_RM_11501_out0 = v_S_9061_out0;
assign v_RM_11503_out0 = v_S_9063_out0;
assign v_RM_11505_out0 = v_S_9065_out0;
assign v_RM_11507_out0 = v_S_9067_out0;
assign v_RM_11509_out0 = v_S_9069_out0;
assign v_RM_11511_out0 = v_S_9071_out0;
assign v_RM_11513_out0 = v_S_9073_out0;
assign v_RM_11515_out0 = v_S_9075_out0;
assign v_RM_11517_out0 = v_S_9077_out0;
assign v_RM_11952_out0 = v_S_9512_out0;
assign v_RM_11954_out0 = v_S_9514_out0;
assign v_RM_11958_out0 = v_S_9518_out0;
assign v_RM_11960_out0 = v_S_9520_out0;
assign v_RM_11962_out0 = v_S_9522_out0;
assign v_RM_11965_out0 = v_S_9525_out0;
assign v_RM_11967_out0 = v_S_9527_out0;
assign v_RM_11969_out0 = v_S_9529_out0;
assign v_RM_11971_out0 = v_S_9531_out0;
assign v_RM_11973_out0 = v_S_9533_out0;
assign v_RM_11975_out0 = v_S_9535_out0;
assign v_RM_11977_out0 = v_S_9537_out0;
assign v_RM_11979_out0 = v_S_9539_out0;
assign v_RM_11981_out0 = v_S_9541_out0;
assign v_MUX1_2717_out0 = v_EXEC2_3241_out0 ? v_REG1_13338_out0 : v__403_out0;
assign v_MUX1_2718_out0 = v_EXEC2_3242_out0 ? v_REG1_13339_out0 : v__404_out0;
assign v_G1_7920_out0 = ((v_RD_6065_out0 && !v_RM_11505_out0) || (!v_RD_6065_out0) && v_RM_11505_out0);
assign v_G1_8384_out0 = ((v_RD_6529_out0 && !v_RM_11969_out0) || (!v_RD_6529_out0) && v_RM_11969_out0);
assign v_G2_12456_out0 = v_RD_6065_out0 && v_RM_11505_out0;
assign v_G2_12920_out0 = v_RD_6529_out0 && v_RM_11969_out0;
assign v_M_REGIN_271_out0 = v_MUX1_2717_out0;
assign v_M_REGIN_272_out0 = v_MUX1_2718_out0;
assign v_CARRY_5065_out0 = v_G2_12456_out0;
assign v_CARRY_5529_out0 = v_G2_12920_out0;
assign v_S_9066_out0 = v_G1_7920_out0;
assign v_S_9530_out0 = v_G1_8384_out0;
assign v_S_1316_out0 = v_S_9066_out0;
assign v_S_1540_out0 = v_S_9530_out0;
assign v_MULTI_REGIN_2870_out0 = v_M_REGIN_271_out0;
assign v_MULTI_REGIN_2871_out0 = v_M_REGIN_272_out0;
assign v_G1_4092_out0 = v_CARRY_5065_out0 || v_CARRY_5064_out0;
assign v_G1_4316_out0 = v_CARRY_5529_out0 || v_CARRY_5528_out0;
assign v_COUT_784_out0 = v_G1_4092_out0;
assign v_COUT_1008_out0 = v_G1_4316_out0;
assign v_MULTI_OUT_13607_out0 = v_MULTI_REGIN_2870_out0;
assign v_MULTI_OUT_13608_out0 = v_MULTI_REGIN_2871_out0;
assign v_MULTI_OUT_1669_out0 = v_MULTI_OUT_13607_out0;
assign v_MULTI_OUT_1670_out0 = v_MULTI_OUT_13608_out0;
assign v_CIN_9911_out0 = v_COUT_784_out0;
assign v_CIN_10135_out0 = v_COUT_1008_out0;
assign v_RD_6077_out0 = v_CIN_9911_out0;
assign v_RD_6541_out0 = v_CIN_10135_out0;
assign v_G1_7932_out0 = ((v_RD_6077_out0 && !v_RM_11517_out0) || (!v_RD_6077_out0) && v_RM_11517_out0);
assign v_G1_8396_out0 = ((v_RD_6541_out0 && !v_RM_11981_out0) || (!v_RD_6541_out0) && v_RM_11981_out0);
assign v_G2_12468_out0 = v_RD_6077_out0 && v_RM_11517_out0;
assign v_G2_12932_out0 = v_RD_6541_out0 && v_RM_11981_out0;
assign v_CARRY_5077_out0 = v_G2_12468_out0;
assign v_CARRY_5541_out0 = v_G2_12932_out0;
assign v_S_9078_out0 = v_G1_7932_out0;
assign v_S_9542_out0 = v_G1_8396_out0;
assign v_S_1322_out0 = v_S_9078_out0;
assign v_S_1546_out0 = v_S_9542_out0;
assign v_G1_4098_out0 = v_CARRY_5077_out0 || v_CARRY_5076_out0;
assign v_G1_4322_out0 = v_CARRY_5541_out0 || v_CARRY_5540_out0;
assign v_COUT_790_out0 = v_G1_4098_out0;
assign v_COUT_1014_out0 = v_G1_4322_out0;
assign v__4788_out0 = { v_S_1316_out0,v_S_1322_out0 };
assign v__4803_out0 = { v_S_1540_out0,v_S_1546_out0 };
assign v_CIN_9906_out0 = v_COUT_790_out0;
assign v_CIN_10130_out0 = v_COUT_1014_out0;
assign v_RD_6067_out0 = v_CIN_9906_out0;
assign v_RD_6531_out0 = v_CIN_10130_out0;
assign v_G1_7922_out0 = ((v_RD_6067_out0 && !v_RM_11507_out0) || (!v_RD_6067_out0) && v_RM_11507_out0);
assign v_G1_8386_out0 = ((v_RD_6531_out0 && !v_RM_11971_out0) || (!v_RD_6531_out0) && v_RM_11971_out0);
assign v_G2_12458_out0 = v_RD_6067_out0 && v_RM_11507_out0;
assign v_G2_12922_out0 = v_RD_6531_out0 && v_RM_11971_out0;
assign v_CARRY_5067_out0 = v_G2_12458_out0;
assign v_CARRY_5531_out0 = v_G2_12922_out0;
assign v_S_9068_out0 = v_G1_7922_out0;
assign v_S_9532_out0 = v_G1_8386_out0;
assign v_S_1317_out0 = v_S_9068_out0;
assign v_S_1541_out0 = v_S_9532_out0;
assign v_G1_4093_out0 = v_CARRY_5067_out0 || v_CARRY_5066_out0;
assign v_G1_4317_out0 = v_CARRY_5531_out0 || v_CARRY_5530_out0;
assign v_COUT_785_out0 = v_G1_4093_out0;
assign v_COUT_1009_out0 = v_G1_4317_out0;
assign v__2558_out0 = { v__4788_out0,v_S_1317_out0 };
assign v__2573_out0 = { v__4803_out0,v_S_1541_out0 };
assign v_CIN_9901_out0 = v_COUT_785_out0;
assign v_CIN_10125_out0 = v_COUT_1009_out0;
assign v_RD_6056_out0 = v_CIN_9901_out0;
assign v_RD_6520_out0 = v_CIN_10125_out0;
assign v_G1_7911_out0 = ((v_RD_6056_out0 && !v_RM_11496_out0) || (!v_RD_6056_out0) && v_RM_11496_out0);
assign v_G1_8375_out0 = ((v_RD_6520_out0 && !v_RM_11960_out0) || (!v_RD_6520_out0) && v_RM_11960_out0);
assign v_G2_12447_out0 = v_RD_6056_out0 && v_RM_11496_out0;
assign v_G2_12911_out0 = v_RD_6520_out0 && v_RM_11960_out0;
assign v_CARRY_5056_out0 = v_G2_12447_out0;
assign v_CARRY_5520_out0 = v_G2_12911_out0;
assign v_S_9057_out0 = v_G1_7911_out0;
assign v_S_9521_out0 = v_G1_8375_out0;
assign v_S_1312_out0 = v_S_9057_out0;
assign v_S_1536_out0 = v_S_9521_out0;
assign v_G1_4088_out0 = v_CARRY_5056_out0 || v_CARRY_5055_out0;
assign v_G1_4312_out0 = v_CARRY_5520_out0 || v_CARRY_5519_out0;
assign v_COUT_780_out0 = v_G1_4088_out0;
assign v_COUT_1004_out0 = v_G1_4312_out0;
assign v__7038_out0 = { v__2558_out0,v_S_1312_out0 };
assign v__7053_out0 = { v__2573_out0,v_S_1536_out0 };
assign v_CIN_9900_out0 = v_COUT_780_out0;
assign v_CIN_10124_out0 = v_COUT_1004_out0;
assign v_RD_6054_out0 = v_CIN_9900_out0;
assign v_RD_6518_out0 = v_CIN_10124_out0;
assign v_G1_7909_out0 = ((v_RD_6054_out0 && !v_RM_11494_out0) || (!v_RD_6054_out0) && v_RM_11494_out0);
assign v_G1_8373_out0 = ((v_RD_6518_out0 && !v_RM_11958_out0) || (!v_RD_6518_out0) && v_RM_11958_out0);
assign v_G2_12445_out0 = v_RD_6054_out0 && v_RM_11494_out0;
assign v_G2_12909_out0 = v_RD_6518_out0 && v_RM_11958_out0;
assign v_CARRY_5054_out0 = v_G2_12445_out0;
assign v_CARRY_5518_out0 = v_G2_12909_out0;
assign v_S_9055_out0 = v_G1_7909_out0;
assign v_S_9519_out0 = v_G1_8373_out0;
assign v_S_1311_out0 = v_S_9055_out0;
assign v_S_1535_out0 = v_S_9519_out0;
assign v_G1_4087_out0 = v_CARRY_5054_out0 || v_CARRY_5053_out0;
assign v_G1_4311_out0 = v_CARRY_5518_out0 || v_CARRY_5517_out0;
assign v_COUT_779_out0 = v_G1_4087_out0;
assign v_COUT_1003_out0 = v_G1_4311_out0;
assign v__13524_out0 = { v__7038_out0,v_S_1311_out0 };
assign v__13539_out0 = { v__7053_out0,v_S_1535_out0 };
assign v_CIN_9907_out0 = v_COUT_779_out0;
assign v_CIN_10131_out0 = v_COUT_1003_out0;
assign v_RD_6069_out0 = v_CIN_9907_out0;
assign v_RD_6533_out0 = v_CIN_10131_out0;
assign v_G1_7924_out0 = ((v_RD_6069_out0 && !v_RM_11509_out0) || (!v_RD_6069_out0) && v_RM_11509_out0);
assign v_G1_8388_out0 = ((v_RD_6533_out0 && !v_RM_11973_out0) || (!v_RD_6533_out0) && v_RM_11973_out0);
assign v_G2_12460_out0 = v_RD_6069_out0 && v_RM_11509_out0;
assign v_G2_12924_out0 = v_RD_6533_out0 && v_RM_11973_out0;
assign v_CARRY_5069_out0 = v_G2_12460_out0;
assign v_CARRY_5533_out0 = v_G2_12924_out0;
assign v_S_9070_out0 = v_G1_7924_out0;
assign v_S_9534_out0 = v_G1_8388_out0;
assign v_S_1318_out0 = v_S_9070_out0;
assign v_S_1542_out0 = v_S_9534_out0;
assign v_G1_4094_out0 = v_CARRY_5069_out0 || v_CARRY_5068_out0;
assign v_G1_4318_out0 = v_CARRY_5533_out0 || v_CARRY_5532_out0;
assign v_COUT_786_out0 = v_G1_4094_out0;
assign v_COUT_1010_out0 = v_G1_4318_out0;
assign v__3317_out0 = { v__13524_out0,v_S_1318_out0 };
assign v__3332_out0 = { v__13539_out0,v_S_1542_out0 };
assign v_CIN_9908_out0 = v_COUT_786_out0;
assign v_CIN_10132_out0 = v_COUT_1010_out0;
assign v_RD_6071_out0 = v_CIN_9908_out0;
assign v_RD_6535_out0 = v_CIN_10132_out0;
assign v_G1_7926_out0 = ((v_RD_6071_out0 && !v_RM_11511_out0) || (!v_RD_6071_out0) && v_RM_11511_out0);
assign v_G1_8390_out0 = ((v_RD_6535_out0 && !v_RM_11975_out0) || (!v_RD_6535_out0) && v_RM_11975_out0);
assign v_G2_12462_out0 = v_RD_6071_out0 && v_RM_11511_out0;
assign v_G2_12926_out0 = v_RD_6535_out0 && v_RM_11975_out0;
assign v_CARRY_5071_out0 = v_G2_12462_out0;
assign v_CARRY_5535_out0 = v_G2_12926_out0;
assign v_S_9072_out0 = v_G1_7926_out0;
assign v_S_9536_out0 = v_G1_8390_out0;
assign v_S_1319_out0 = v_S_9072_out0;
assign v_S_1543_out0 = v_S_9536_out0;
assign v_G1_4095_out0 = v_CARRY_5071_out0 || v_CARRY_5070_out0;
assign v_G1_4319_out0 = v_CARRY_5535_out0 || v_CARRY_5534_out0;
assign v_COUT_787_out0 = v_G1_4095_out0;
assign v_COUT_1011_out0 = v_G1_4319_out0;
assign v__7153_out0 = { v__3317_out0,v_S_1319_out0 };
assign v__7168_out0 = { v__3332_out0,v_S_1543_out0 };
assign v_CIN_9910_out0 = v_COUT_787_out0;
assign v_CIN_10134_out0 = v_COUT_1011_out0;
assign v_RD_6075_out0 = v_CIN_9910_out0;
assign v_RD_6539_out0 = v_CIN_10134_out0;
assign v_G1_7930_out0 = ((v_RD_6075_out0 && !v_RM_11515_out0) || (!v_RD_6075_out0) && v_RM_11515_out0);
assign v_G1_8394_out0 = ((v_RD_6539_out0 && !v_RM_11979_out0) || (!v_RD_6539_out0) && v_RM_11979_out0);
assign v_G2_12466_out0 = v_RD_6075_out0 && v_RM_11515_out0;
assign v_G2_12930_out0 = v_RD_6539_out0 && v_RM_11979_out0;
assign v_CARRY_5075_out0 = v_G2_12466_out0;
assign v_CARRY_5539_out0 = v_G2_12930_out0;
assign v_S_9076_out0 = v_G1_7930_out0;
assign v_S_9540_out0 = v_G1_8394_out0;
assign v_S_1321_out0 = v_S_9076_out0;
assign v_S_1545_out0 = v_S_9540_out0;
assign v_G1_4097_out0 = v_CARRY_5075_out0 || v_CARRY_5074_out0;
assign v_G1_4321_out0 = v_CARRY_5539_out0 || v_CARRY_5538_out0;
assign v_COUT_789_out0 = v_G1_4097_out0;
assign v_COUT_1013_out0 = v_G1_4321_out0;
assign v__4755_out0 = { v__7153_out0,v_S_1321_out0 };
assign v__4770_out0 = { v__7168_out0,v_S_1545_out0 };
assign v_CIN_9903_out0 = v_COUT_789_out0;
assign v_CIN_10127_out0 = v_COUT_1013_out0;
assign v_RD_6061_out0 = v_CIN_9903_out0;
assign v_RD_6525_out0 = v_CIN_10127_out0;
assign v_G1_7916_out0 = ((v_RD_6061_out0 && !v_RM_11501_out0) || (!v_RD_6061_out0) && v_RM_11501_out0);
assign v_G1_8380_out0 = ((v_RD_6525_out0 && !v_RM_11965_out0) || (!v_RD_6525_out0) && v_RM_11965_out0);
assign v_G2_12452_out0 = v_RD_6061_out0 && v_RM_11501_out0;
assign v_G2_12916_out0 = v_RD_6525_out0 && v_RM_11965_out0;
assign v_CARRY_5061_out0 = v_G2_12452_out0;
assign v_CARRY_5525_out0 = v_G2_12916_out0;
assign v_S_9062_out0 = v_G1_7916_out0;
assign v_S_9526_out0 = v_G1_8380_out0;
assign v_S_1314_out0 = v_S_9062_out0;
assign v_S_1538_out0 = v_S_9526_out0;
assign v_G1_4090_out0 = v_CARRY_5061_out0 || v_CARRY_5060_out0;
assign v_G1_4314_out0 = v_CARRY_5525_out0 || v_CARRY_5524_out0;
assign v_COUT_782_out0 = v_G1_4090_out0;
assign v_COUT_1006_out0 = v_G1_4314_out0;
assign v__6932_out0 = { v__4755_out0,v_S_1314_out0 };
assign v__6947_out0 = { v__4770_out0,v_S_1538_out0 };
assign v_CIN_9904_out0 = v_COUT_782_out0;
assign v_CIN_10128_out0 = v_COUT_1006_out0;
assign v_RD_6063_out0 = v_CIN_9904_out0;
assign v_RD_6527_out0 = v_CIN_10128_out0;
assign v_G1_7918_out0 = ((v_RD_6063_out0 && !v_RM_11503_out0) || (!v_RD_6063_out0) && v_RM_11503_out0);
assign v_G1_8382_out0 = ((v_RD_6527_out0 && !v_RM_11967_out0) || (!v_RD_6527_out0) && v_RM_11967_out0);
assign v_G2_12454_out0 = v_RD_6063_out0 && v_RM_11503_out0;
assign v_G2_12918_out0 = v_RD_6527_out0 && v_RM_11967_out0;
assign v_CARRY_5063_out0 = v_G2_12454_out0;
assign v_CARRY_5527_out0 = v_G2_12918_out0;
assign v_S_9064_out0 = v_G1_7918_out0;
assign v_S_9528_out0 = v_G1_8382_out0;
assign v_S_1315_out0 = v_S_9064_out0;
assign v_S_1539_out0 = v_S_9528_out0;
assign v_G1_4091_out0 = v_CARRY_5063_out0 || v_CARRY_5062_out0;
assign v_G1_4315_out0 = v_CARRY_5527_out0 || v_CARRY_5526_out0;
assign v_COUT_783_out0 = v_G1_4091_out0;
assign v_COUT_1007_out0 = v_G1_4315_out0;
assign v__5808_out0 = { v__6932_out0,v_S_1315_out0 };
assign v__5823_out0 = { v__6947_out0,v_S_1539_out0 };
assign v_CIN_9909_out0 = v_COUT_783_out0;
assign v_CIN_10133_out0 = v_COUT_1007_out0;
assign v_RD_6073_out0 = v_CIN_9909_out0;
assign v_RD_6537_out0 = v_CIN_10133_out0;
assign v_G1_7928_out0 = ((v_RD_6073_out0 && !v_RM_11513_out0) || (!v_RD_6073_out0) && v_RM_11513_out0);
assign v_G1_8392_out0 = ((v_RD_6537_out0 && !v_RM_11977_out0) || (!v_RD_6537_out0) && v_RM_11977_out0);
assign v_G2_12464_out0 = v_RD_6073_out0 && v_RM_11513_out0;
assign v_G2_12928_out0 = v_RD_6537_out0 && v_RM_11977_out0;
assign v_CARRY_5073_out0 = v_G2_12464_out0;
assign v_CARRY_5537_out0 = v_G2_12928_out0;
assign v_S_9074_out0 = v_G1_7928_out0;
assign v_S_9538_out0 = v_G1_8392_out0;
assign v_S_1320_out0 = v_S_9074_out0;
assign v_S_1544_out0 = v_S_9538_out0;
assign v_G1_4096_out0 = v_CARRY_5073_out0 || v_CARRY_5072_out0;
assign v_G1_4320_out0 = v_CARRY_5537_out0 || v_CARRY_5536_out0;
assign v_COUT_788_out0 = v_G1_4096_out0;
assign v_COUT_1012_out0 = v_G1_4320_out0;
assign v__2032_out0 = { v__5808_out0,v_S_1320_out0 };
assign v__2047_out0 = { v__5823_out0,v_S_1544_out0 };
assign v_CIN_9897_out0 = v_COUT_788_out0;
assign v_CIN_10121_out0 = v_COUT_1012_out0;
assign v_RD_6048_out0 = v_CIN_9897_out0;
assign v_RD_6512_out0 = v_CIN_10121_out0;
assign v_G1_7903_out0 = ((v_RD_6048_out0 && !v_RM_11488_out0) || (!v_RD_6048_out0) && v_RM_11488_out0);
assign v_G1_8367_out0 = ((v_RD_6512_out0 && !v_RM_11952_out0) || (!v_RD_6512_out0) && v_RM_11952_out0);
assign v_G2_12439_out0 = v_RD_6048_out0 && v_RM_11488_out0;
assign v_G2_12903_out0 = v_RD_6512_out0 && v_RM_11952_out0;
assign v_CARRY_5048_out0 = v_G2_12439_out0;
assign v_CARRY_5512_out0 = v_G2_12903_out0;
assign v_S_9049_out0 = v_G1_7903_out0;
assign v_S_9513_out0 = v_G1_8367_out0;
assign v_S_1308_out0 = v_S_9049_out0;
assign v_S_1532_out0 = v_S_9513_out0;
assign v_G1_4084_out0 = v_CARRY_5048_out0 || v_CARRY_5047_out0;
assign v_G1_4308_out0 = v_CARRY_5512_out0 || v_CARRY_5511_out0;
assign v_COUT_776_out0 = v_G1_4084_out0;
assign v_COUT_1000_out0 = v_G1_4308_out0;
assign v__2799_out0 = { v__2032_out0,v_S_1308_out0 };
assign v__2814_out0 = { v__2047_out0,v_S_1532_out0 };
assign v_CIN_9902_out0 = v_COUT_776_out0;
assign v_CIN_10126_out0 = v_COUT_1000_out0;
assign v_RD_6058_out0 = v_CIN_9902_out0;
assign v_RD_6522_out0 = v_CIN_10126_out0;
assign v_G1_7913_out0 = ((v_RD_6058_out0 && !v_RM_11498_out0) || (!v_RD_6058_out0) && v_RM_11498_out0);
assign v_G1_8377_out0 = ((v_RD_6522_out0 && !v_RM_11962_out0) || (!v_RD_6522_out0) && v_RM_11962_out0);
assign v_G2_12449_out0 = v_RD_6058_out0 && v_RM_11498_out0;
assign v_G2_12913_out0 = v_RD_6522_out0 && v_RM_11962_out0;
assign v_CARRY_5058_out0 = v_G2_12449_out0;
assign v_CARRY_5522_out0 = v_G2_12913_out0;
assign v_S_9059_out0 = v_G1_7913_out0;
assign v_S_9523_out0 = v_G1_8377_out0;
assign v_S_1313_out0 = v_S_9059_out0;
assign v_S_1537_out0 = v_S_9523_out0;
assign v_G1_4089_out0 = v_CARRY_5058_out0 || v_CARRY_5057_out0;
assign v_G1_4313_out0 = v_CARRY_5522_out0 || v_CARRY_5521_out0;
assign v_COUT_781_out0 = v_G1_4089_out0;
assign v_COUT_1005_out0 = v_G1_4313_out0;
assign v__1831_out0 = { v__2799_out0,v_S_1313_out0 };
assign v__1846_out0 = { v__2814_out0,v_S_1537_out0 };
assign v_CIN_9898_out0 = v_COUT_781_out0;
assign v_CIN_10122_out0 = v_COUT_1005_out0;
assign v_RD_6050_out0 = v_CIN_9898_out0;
assign v_RD_6514_out0 = v_CIN_10122_out0;
assign v_G1_7905_out0 = ((v_RD_6050_out0 && !v_RM_11490_out0) || (!v_RD_6050_out0) && v_RM_11490_out0);
assign v_G1_8369_out0 = ((v_RD_6514_out0 && !v_RM_11954_out0) || (!v_RD_6514_out0) && v_RM_11954_out0);
assign v_G2_12441_out0 = v_RD_6050_out0 && v_RM_11490_out0;
assign v_G2_12905_out0 = v_RD_6514_out0 && v_RM_11954_out0;
assign v_CARRY_5050_out0 = v_G2_12441_out0;
assign v_CARRY_5514_out0 = v_G2_12905_out0;
assign v_S_9051_out0 = v_G1_7905_out0;
assign v_S_9515_out0 = v_G1_8369_out0;
assign v_S_1309_out0 = v_S_9051_out0;
assign v_S_1533_out0 = v_S_9515_out0;
assign v_G1_4085_out0 = v_CARRY_5050_out0 || v_CARRY_5049_out0;
assign v_G1_4309_out0 = v_CARRY_5514_out0 || v_CARRY_5513_out0;
assign v_COUT_777_out0 = v_G1_4085_out0;
assign v_COUT_1001_out0 = v_G1_4309_out0;
assign v__4555_out0 = { v__1831_out0,v_S_1309_out0 };
assign v__4570_out0 = { v__1846_out0,v_S_1533_out0 };
assign v_RM_3446_out0 = v_COUT_777_out0;
assign v_RM_3670_out0 = v_COUT_1001_out0;
assign v_RM_11491_out0 = v_RM_3446_out0;
assign v_RM_11955_out0 = v_RM_3670_out0;
assign v_G1_7906_out0 = ((v_RD_6051_out0 && !v_RM_11491_out0) || (!v_RD_6051_out0) && v_RM_11491_out0);
assign v_G1_8370_out0 = ((v_RD_6515_out0 && !v_RM_11955_out0) || (!v_RD_6515_out0) && v_RM_11955_out0);
assign v_G2_12442_out0 = v_RD_6051_out0 && v_RM_11491_out0;
assign v_G2_12906_out0 = v_RD_6515_out0 && v_RM_11955_out0;
assign v_CARRY_5051_out0 = v_G2_12442_out0;
assign v_CARRY_5515_out0 = v_G2_12906_out0;
assign v_S_9052_out0 = v_G1_7906_out0;
assign v_S_9516_out0 = v_G1_8370_out0;
assign v_RM_11492_out0 = v_S_9052_out0;
assign v_RM_11956_out0 = v_S_9516_out0;
assign v_G1_7907_out0 = ((v_RD_6052_out0 && !v_RM_11492_out0) || (!v_RD_6052_out0) && v_RM_11492_out0);
assign v_G1_8371_out0 = ((v_RD_6516_out0 && !v_RM_11956_out0) || (!v_RD_6516_out0) && v_RM_11956_out0);
assign v_G2_12443_out0 = v_RD_6052_out0 && v_RM_11492_out0;
assign v_G2_12907_out0 = v_RD_6516_out0 && v_RM_11956_out0;
assign v_CARRY_5052_out0 = v_G2_12443_out0;
assign v_CARRY_5516_out0 = v_G2_12907_out0;
assign v_S_9053_out0 = v_G1_7907_out0;
assign v_S_9517_out0 = v_G1_8371_out0;
assign v_S_1310_out0 = v_S_9053_out0;
assign v_S_1534_out0 = v_S_9517_out0;
assign v_G1_4086_out0 = v_CARRY_5052_out0 || v_CARRY_5051_out0;
assign v_G1_4310_out0 = v_CARRY_5516_out0 || v_CARRY_5515_out0;
assign v_COUT_778_out0 = v_G1_4086_out0;
assign v_COUT_1002_out0 = v_G1_4310_out0;
assign v__10657_out0 = { v__4555_out0,v_S_1310_out0 };
assign v__10672_out0 = { v__4570_out0,v_S_1534_out0 };
assign v__10952_out0 = { v__10657_out0,v_COUT_778_out0 };
assign v__10967_out0 = { v__10672_out0,v_COUT_1002_out0 };
assign v_COUT_10922_out0 = v__10952_out0;
assign v_COUT_10937_out0 = v__10967_out0;
assign v__212_out0 = { v__403_out0,v_COUT_10922_out0 };
assign v__213_out0 = { v__404_out0,v_COUT_10937_out0 };
assign v_FLOATING_MULTI_7697_out0 = v__212_out0;
assign v_FLOATING_MULTI_7698_out0 = v__213_out0;
assign v_32BIT_MULTI_1183_out0 = v_FLOATING_MULTI_7697_out0;
assign v_32BIT_MULTI_1184_out0 = v_FLOATING_MULTI_7698_out0;
assign v_32BITPRODUCT_82_out0 = v_32BIT_MULTI_1183_out0;
assign v_32BITPRODUCT_83_out0 = v_32BIT_MULTI_1184_out0;
assign v_32BITPRODUCT_12249_out0 = v_32BITPRODUCT_82_out0;
assign v_32BITPRODUCT_12250_out0 = v_32BITPRODUCT_83_out0;
assign v_SEL7_4850_out0 = v_32BITPRODUCT_12249_out0[21:10];
assign v_SEL7_4851_out0 = v_32BITPRODUCT_12250_out0[21:10];
assign v_MULTI_PRODUCT_7104_out0 = v_SEL7_4850_out0;
assign v_MULTI_PRODUCT_7105_out0 = v_SEL7_4851_out0;
assign v_MUX8_13785_out0 = v_MULTI_INSTRUCTION_2451_out0 ? v_MULTI_PRODUCT_7104_out0 : v_SEL8_10686_out0;
assign v_MUX8_13786_out0 = v_MULTI_INSTRUCTION_2452_out0 ? v_MULTI_PRODUCT_7105_out0 : v_SEL8_10687_out0;
assign v_SEL3_1143_out0 = v_MUX8_13785_out0[11:11];
assign v_SEL3_1144_out0 = v_MUX8_13786_out0[11:11];
assign v_SEL5_3049_out0 = v_MUX8_13785_out0[10:10];
assign v_SEL5_3050_out0 = v_MUX8_13786_out0[10:10];
assign v_SEL2_13496_out0 = v_MUX8_13785_out0[10:0];
assign v_SEL2_13497_out0 = v_MUX8_13786_out0[10:0];
assign v_SEL6_3991_out0 = v_SEL2_13496_out0[8:0];
assign v_SEL6_3992_out0 = v_SEL2_13497_out0[8:0];
assign v_BIT10_7009_out0 = v_SEL5_3049_out0;
assign v_BIT10_7010_out0 = v_SEL5_3050_out0;
assign v_OVERFLOW_10492_out0 = v_SEL3_1143_out0;
assign v_OVERFLOW_10493_out0 = v_SEL3_1144_out0;
assign v_SEL4_11225_out0 = v_SEL2_13496_out0[9:0];
assign v_SEL4_11226_out0 = v_SEL2_13497_out0[9:0];
assign v_SEL9_13753_out0 = v_SEL2_13496_out0[10:1];
assign v_SEL9_13754_out0 = v_SEL2_13497_out0[10:1];
assign v_G3_2690_out0 = v_BIT10_7009_out0 || v_OVERFLOW_10492_out0;
assign v_G3_2691_out0 = v_BIT10_7010_out0 || v_OVERFLOW_10493_out0;
assign v__8677_out0 = { v_C9_3029_out0,v_SEL6_3991_out0 };
assign v__8678_out0 = { v_C9_3030_out0,v_SEL6_3992_out0 };
assign v_MUX5_10260_out0 = v_SUBNORMAL_8808_out0 ? v_BIT10_7009_out0 : v_OVERFLOW_10492_out0;
assign v_MUX5_10261_out0 = v_SUBNORMAL_8809_out0 ? v_BIT10_7010_out0 : v_OVERFLOW_10493_out0;
assign v_MUX4_10357_out0 = v_OVERFLOW_10492_out0 ? v_SEL9_13753_out0 : v_SEL4_11225_out0;
assign v_MUX4_10358_out0 = v_OVERFLOW_10493_out0 ? v_SEL9_13754_out0 : v_SEL4_11226_out0;
assign v_G2_5840_out0 = !(v_G3_2690_out0 || v_SUBNORMAL_8808_out0);
assign v_G2_5841_out0 = !(v_G3_2691_out0 || v_SUBNORMAL_8809_out0);
assign v_UNDERFLOW_6916_out0 = v_G2_5840_out0;
assign v_UNDERFLOW_6917_out0 = v_G2_5841_out0;
assign v_G4_3235_out0 = v_UNDERFLOW_6916_out0 && v_G5_638_out0;
assign v_G4_3236_out0 = v_UNDERFLOW_6917_out0 && v_G5_639_out0;
assign v_MUX7_4481_out0 = v_UNDERFLOW_6916_out0 ? v_C10_11248_out0 : v_C8_2758_out0;
assign v_MUX7_4482_out0 = v_UNDERFLOW_6917_out0 ? v_C10_11249_out0 : v_C8_2759_out0;
assign {v_A7_2719_out1,v_A7_2719_out0 } = v_EXP_2441_out0 + v_MUX7_4481_out0 + v_MUX5_10260_out0;
assign {v_A7_2720_out1,v_A7_2720_out0 } = v_EXP_2442_out0 + v_MUX7_4482_out0 + v_MUX5_10261_out0;
assign v_MUX6_10350_out0 = v_G4_3235_out0 ? v__8677_out0 : v_MUX4_10357_out0;
assign v_MUX6_10351_out0 = v_G4_3236_out0 ? v__8678_out0 : v_MUX4_10358_out0;
assign v_SIG_ANS_439_out0 = v_MUX6_10350_out0;
assign v_SIG_ANS_440_out0 = v_MUX6_10351_out0;
assign v_NOTUSED3_10550_out0 = v_A7_2719_out1;
assign v_NOTUSED3_10551_out0 = v_A7_2720_out1;
assign v_EXP_ANS_13748_out0 = v_A7_2719_out0;
assign v_EXP_ANS_13749_out0 = v_A7_2720_out0;
assign v_EXP_ANS_2008_out0 = v_EXP_ANS_13748_out0;
assign v_EXP_ANS_2009_out0 = v_EXP_ANS_13749_out0;
assign v_SIG_ANS_2335_out0 = v_SIG_ANS_439_out0;
assign v_SIG_ANS_2336_out0 = v_SIG_ANS_440_out0;
assign v__2610_out0 = { v_EXP_ANS_2008_out0,v_SIGN_ANS_8650_out0 };
assign v__2611_out0 = { v_EXP_ANS_2009_out0,v_SIGN_ANS_8651_out0 };
assign v_SIG_ANS_3276_out0 = v_SIG_ANS_2335_out0;
assign v_SIG_ANS_3277_out0 = v_SIG_ANS_2336_out0;
assign v_EXP_ANS_10487_out0 = v_EXP_ANS_2008_out0;
assign v_EXP_ANS_10488_out0 = v_EXP_ANS_2009_out0;
assign v_SIG_ANS_10296_out0 = v_SIG_ANS_3276_out0;
assign v_SIG_ANS_10297_out0 = v_SIG_ANS_3277_out0;
assign v__10449_out0 = { v_SIG_ANS_2335_out0,v__2610_out0 };
assign v__10450_out0 = { v_SIG_ANS_2336_out0,v__2611_out0 };
assign v_EXP_ANS_11059_out0 = v_EXP_ANS_10487_out0;
assign v_EXP_ANS_11060_out0 = v_EXP_ANS_10488_out0;
assign v_16BIT_WORD_ANSWER_8821_out0 = v__10449_out0;
assign v_16BIT_WORD_ANSWER_8822_out0 = v__10450_out0;
assign v_FLOATING_REGISTER_IN_562_out0 = v_16BIT_WORD_ANSWER_8821_out0;
assign v_FLOATING_REGISTER_IN_563_out0 = v_16BIT_WORD_ANSWER_8822_out0;
assign v_MUX12_1714_out0 = v_FLOATING_EN_ALU_634_out0 ? v_FLOATING_REGISTER_IN_562_out0 : v_ALUOUT_4607_out0;
assign v_MUX12_1715_out0 = v_FLOATING_EN_ALU_635_out0 ? v_FLOATING_REGISTER_IN_563_out0 : v_ALUOUT_4608_out0;
assign v_MUX5_2606_out0 = v_FLOATING_INS_13797_out0 ? v_FLOATING_REGISTER_IN_562_out0 : v_MULTI_REGIN_2870_out0;
assign v_MUX5_2607_out0 = v_FLOATING_INS_13798_out0 ? v_FLOATING_REGISTER_IN_563_out0 : v_MULTI_REGIN_2871_out0;
assign v_MUX4_10_out0 = v_MULTI_OPCODE_3020_out0 ? v_MUX5_2606_out0 : v_LS_REGIN_3303_out0;
assign v_MUX4_11_out0 = v_MULTI_OPCODE_3021_out0 ? v_MUX5_2607_out0 : v_LS_REGIN_3304_out0;
assign v_MUX11_13745_out0 = v_IR15_2464_out0 ? v_MUX12_1714_out0 : v_MUX4_10_out0;
assign v_MUX11_13746_out0 = v_IR15_2465_out0 ? v_MUX12_1715_out0 : v_MUX4_11_out0;
assign v_DIN_2266_out0 = v_MUX11_13745_out0;
assign v_DIN_2267_out0 = v_MUX11_13746_out0;
assign v_DIN3_10310_out0 = v_MUX11_13745_out0;
assign v_DIN3_10311_out0 = v_MUX11_13746_out0;
assign v_DIN_9798_out0 = v_DIN_2266_out0;
assign v_DIN_9799_out0 = v_DIN_2267_out0;


endmodule
